CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 370 30 80 10
2 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
170 176 283 273
9437202 0
0
6 Title:
5 Name:
0
0
0
72
13 Logic Switch~
5 923 1458 0 10 11
0 11 0 0 0 0 0 0 0 0
1
0
0 0 21360 692
2 5V
-7 -16 7 -8
3 V13
-11 -26 10 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7670 0 0
2
43336.5 0
0
13 Logic Switch~
5 961 1373 0 1 11
0 40
0
0 0 21360 90
2 0V
9 0 23 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
951 0 0
2
43336.5 1
0
13 Logic Switch~
5 913 1372 0 1 11
0 41
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9536 0 0
2
43336.5 2
0
13 Logic Switch~
5 549 154 0 1 11
0 55
0
0 0 21360 0
2 0V
-8 -17 6 -9
3 V11
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5495 0 0
2
43336.5 3
0
13 Logic Switch~
5 550 669 0 1 11
0 16
0
0 0 21360 0
2 0V
-8 -16 6 -8
3 V10
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8152 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 553 597 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6223 0 0
2
5.89859e-315 5.26354e-315
0
13 Logic Switch~
5 554 536 0 1 11
0 20
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V8
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5441 0 0
2
5.89859e-315 5.30499e-315
0
13 Logic Switch~
5 551 480 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3189 0 0
2
5.89859e-315 5.32571e-315
0
13 Logic Switch~
5 553 401 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8460 0 0
2
5.89859e-315 5.34643e-315
0
13 Logic Switch~
5 551 342 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5179 0 0
2
5.89859e-315 5.3568e-315
0
13 Logic Switch~
5 552 269 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3593 0 0
2
5.89859e-315 5.36716e-315
0
13 Logic Switch~
5 551 214 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -19 7 -11
2 V3
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3928 0 0
2
5.89859e-315 5.37752e-315
0
7 Ground~
168 1163 1085 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
363 0 0
2
43336.5 0
0
7 74LS157
122 1202 1017 0 14 29
0 11 15 10 14 9 13 8 12 7
2 6 5 4 3
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
3 U18
-11 -61 10 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
8132 0 0
2
43336.5 0
0
14 Logic Display~
6 1287 1160 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
65 0 0
2
43336.5 4
0
14 Logic Display~
6 1285 1088 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6609 0 0
2
43336.5 5
0
14 Logic Display~
6 1284 1031 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8995 0 0
2
43336.5 6
0
14 Logic Display~
6 1284 975 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3918 0 0
2
43336.5 7
0
14 Logic Display~
6 984 1292 0 1 2
10 12
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7519 0 0
2
43336.5 16
0
14 Logic Display~
6 980 1137 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
377 0 0
2
43336.5 17
0
14 Logic Display~
6 979 1003 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8816 0 0
2
43336.5 18
0
14 Logic Display~
6 975 870 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3877 0 0
2
43336.5 19
0
5 4049~
219 694 1192 0 2 22
0 17 33
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
926 0 0
2
43336.5 20
0
5 4049~
219 683 1046 0 2 22
0 19 30
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
7262 0 0
2
43336.5 21
0
5 4049~
219 675 760 0 2 22
0 23 24
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 1 0
1 U
5267 0 0
2
43336.5 22
0
5 4049~
219 679 905 0 2 22
0 21 27
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 1 0
1 U
8838 0 0
2
43336.5 23
0
5 4081~
219 780 1270 0 3 22
0 17 16 35
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
7159 0 0
2
43336.5 24
0
5 4081~
219 768 1118 0 3 22
0 19 18 32
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
5812 0 0
2
43336.5 25
0
5 4081~
219 750 837 0 3 22
0 23 22 26
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
331 0 0
2
43336.5 26
0
5 4081~
219 758 978 0 3 22
0 21 20 29
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U16A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
9604 0 0
2
43336.5 27
0
5 4030~
219 692 1232 0 3 22
0 17 16 34
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U15D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
7518 0 0
2
43336.5 28
0
5 4030~
219 684 1086 0 3 22
0 19 18 31
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U15C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
4832 0 0
2
43336.5 29
0
5 4030~
219 678 949 0 3 22
0 21 20 28
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U15B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
6798 0 0
2
43336.5 30
0
5 4030~
219 676 802 0 3 22
0 23 22 25
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U15A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3336 0 0
2
43336.5 31
0
5 4071~
219 766 1320 0 3 22
0 17 16 36
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11D
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
8370 0 0
2
43336.5 32
0
5 4071~
219 760 1166 0 3 22
0 19 18 37
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3910 0 0
2
43336.5 33
0
5 4071~
219 752 1026 0 3 22
0 21 20 38
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
316 0 0
2
43336.5 34
0
7 74LS151
20 856 1281 0 14 29
0 56 57 58 59 33 34 35 36 2
2 41 40 12 60
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U14
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
536 0 0
2
43336.5 35
0
7 Ground~
168 954 1264 0 1 3
0 2
0
0 0 53360 0
0
5 GND10
-17 -26 18 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4460 0 0
2
43336.5 36
0
7 74LS151
20 852 1130 0 14 29
0 61 62 63 64 30 31 32 37 2
2 41 40 13 65
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3260 0 0
2
43336.5 37
0
7 Ground~
168 952 1112 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5156 0 0
2
43336.5 38
0
7 74LS151
20 851 990 0 14 29
0 66 67 68 69 27 28 29 38 2
2 41 40 14 70
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U12
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3133 0 0
2
43336.5 39
0
7 Ground~
168 949 973 0 1 3
0 2
0
0 0 53360 0
0
4 GND8
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5523 0 0
2
43336.5 40
0
5 4071~
219 744 886 0 3 22
0 23 22 39
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U11A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
3746 0 0
2
43336.5 41
0
7 Ground~
168 945 839 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5668 0 0
2
43336.5 42
0
7 74LS151
20 847 850 0 14 29
0 71 72 73 74 24 25 26 39 2
2 41 40 15 75
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U10
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
5368 0 0
2
43336.5 43
0
14 Logic Display~
6 1135 658 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8293 0 0
2
43336.5 44
0
7 Ground~
168 945 653 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3232 0 0
2
43336.5 45
0
7 Ground~
168 898 510 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6644 0 0
2
43336.5 46
0
7 Ground~
168 894 385 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
4978 0 0
2
43336.5 47
0
7 Ground~
168 897 236 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9207 0 0
2
43336.5 48
0
7 74LS151
20 840 669 0 14 29
0 76 77 78 79 46 50 16 2 2
2 41 40 42 80
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
6998 0 0
2
43336.5 49
0
7 74LS151
20 836 528 0 14 29
0 81 82 83 84 46 49 18 2 2
2 41 40 43 85
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U7
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3175 0 0
2
43336.5 50
0
7 74LS151
20 832 402 0 14 29
0 86 87 88 89 46 48 20 2 2
2 41 40 44 90
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U6
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3378 0 0
2
43336.5 51
0
7 74LS151
20 830 248 0 14 29
0 91 92 93 94 46 47 22 2 2
2 41 40 45 95
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
2 U5
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
922 0 0
2
43336.5 52
0
5 4049~
219 691 669 0 2 22
0 16 50
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 1 0
1 U
6891 0 0
2
43336.5 53
0
5 4049~
219 695 518 0 2 22
0 18 49
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 1 0
1 U
5407 0 0
2
43336.5 54
0
5 4049~
219 689 406 0 2 22
0 20 48
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 1 0
1 U
7349 0 0
2
43336.5 55
0
5 4049~
219 684 244 0 2 22
0 22 47
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U9A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 1 0
1 U
3919 0 0
2
43336.5 56
0
7 Ground~
168 769 120 0 1 3
0 2
0
0 0 53360 180
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9747 0 0
2
43336.5 57
0
8 Battery~
219 728 120 0 2 5
0 96 46
0
0 0 880 0
2 5V
15 -2 29 6
3 V12
11 -15 32 -7
0
0
14 %D %1 %2 DC %V
0
0
0
5

0 1 2 1 2 0
86 0 0 512 1 0 0 0
1 V
5310 0 0
2
43336.5 58
0
12 Hex Display~
7 1178 484 0 18 19
10 10 9 8 7 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4318 0 0
2
43336.5 59
0
14 Logic Display~
6 1137 729 0 1 2
10 51
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3917 0 0
2
43336.5 60
0
12 Hex Display~
7 428 484 0 16 19
10 22 20 18 16 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7930 0 0
2
43336.5 61
0
12 Hex Display~
7 447 203 0 18 19
10 23 21 19 17 0 0 0 0 0
0 0 1 1 0 0 0 0 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
6128 0 0
2
43336.5 62
0
14 Logic Display~
6 1125 491 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7346 0 0
2
43336.5 63
0
14 Logic Display~
6 1123 346 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8577 0 0
2
43336.5 64
0
14 Logic Display~
6 1121 178 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3372 0 0
2
43336.5 65
0
4 4008
219 1033 240 0 14 29
0 97 98 99 23 100 101 102 45 55
10 54 103 104 105
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3741 0 0
2
5.89859e-315 5.38788e-315
0
4 4008
219 1034 369 0 14 29
0 106 107 108 21 109 110 111 44 54
9 53 112 113 114
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
5813 0 0
2
5.89859e-315 5.39306e-315
0
4 4008
219 1032 510 0 14 29
0 115 116 117 19 118 119 120 43 53
8 52 121 122 123
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3213 0 0
2
5.89859e-315 5.39824e-315
0
4 4008
219 1033 680 0 14 29
0 124 125 126 17 127 128 129 42 52
7 51 130 131 132
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3694 0 0
2
5.89859e-315 5.40342e-315
0
144
1 10 2 0 0 12288 0 13 14 0 0 5
1163 1079
1163 1073
1162 1073
1162 1062
1164 1062
14 1 3 0 0 8320 0 14 15 0 0 5
1234 1053
1262 1053
1262 1206
1287 1206
1287 1178
13 1 4 0 0 8320 0 14 16 0 0 5
1234 1035
1267 1035
1267 1134
1285 1134
1285 1106
12 1 5 0 0 8320 0 14 17 0 0 5
1234 1017
1271 1017
1271 1057
1284 1057
1284 1049
11 1 6 0 0 4224 0 14 18 0 0 3
1234 999
1284 999
1284 993
0 9 7 0 0 4240 0 0 14 126 0 3
1125 689
1125 1053
1170 1053
0 7 8 0 0 4224 0 0 14 82 0 3
1150 519
1150 1035
1170 1035
0 5 9 0 0 4224 0 0 14 127 0 3
1162 513
1162 1017
1170 1017
0 3 10 0 0 4224 0 0 14 128 0 5
1195 508
1195 959
1153 959
1153 999
1170 999
1 1 11 0 0 8320 0 1 14 0 0 4
935 1458
1143 1458
1143 981
1170 981
1 8 12 0 0 12416 0 19 14 0 0 5
984 1310
984 1319
1153 1319
1153 1044
1170 1044
0 6 13 0 0 4224 0 0 14 16 0 4
980 1159
1148 1159
1148 1026
1170 1026
1 4 14 0 0 8320 0 21 14 0 0 5
979 1021
979 1028
1153 1028
1153 1008
1170 1008
0 2 15 0 0 8320 0 0 14 18 0 3
974 896
974 990
1170 990
1 13 12 0 0 0 0 19 38 0 0 5
984 1310
984 1314
902 1314
902 1308
888 1308
1 13 13 0 0 0 0 20 40 0 0 5
980 1155
980 1159
898 1159
898 1157
884 1157
1 13 14 0 0 0 0 21 42 0 0 5
979 1021
979 1025
897 1025
897 1017
883 1017
13 1 15 0 0 0 0 46 22 0 0 5
879 877
963 877
963 896
975 896
975 888
0 2 16 0 0 12288 0 0 35 20 0 4
642 1284
643 1284
643 1329
753 1329
0 2 16 0 0 16384 0 0 27 21 0 5
642 1241
642 1284
642 1284
642 1279
756 1279
0 2 16 0 0 4224 0 0 31 133 0 3
567 669
567 1241
676 1241
0 1 17 0 0 12288 0 0 35 23 0 4
659 1267
658 1267
658 1311
753 1311
0 1 17 0 0 20480 0 0 27 24 0 6
660 1221
659 1221
659 1267
659 1267
659 1261
756 1261
0 1 17 0 0 0 0 0 31 43 0 3
660 1192
660 1223
676 1223
0 2 18 0 0 4096 0 0 36 26 0 3
729 1127
729 1175
747 1175
2 0 18 0 0 4096 0 28 0 0 40 3
744 1127
654 1127
654 1095
0 1 19 0 0 4096 0 0 36 28 0 3
719 1109
719 1157
747 1157
0 1 19 0 0 12288 0 0 28 29 0 4
647 1076
650 1076
650 1109
744 1109
0 1 19 0 0 0 0 0 32 44 0 3
647 1046
647 1077
668 1077
0 2 20 0 0 4096 0 0 37 31 0 5
691 987
691 1032
731 1032
731 1035
739 1035
0 2 20 0 0 8192 0 0 30 41 0 3
643 958
643 987
734 987
0 1 21 0 0 4096 0 0 37 33 0 3
700 969
700 1017
739 1017
0 1 21 0 0 12288 0 0 30 34 0 4
640 940
658 940
658 969
734 969
0 1 21 0 0 0 0 0 33 45 0 3
640 905
640 940
662 940
0 2 22 0 0 4096 0 0 44 36 0 3
709 846
709 895
731 895
0 2 22 0 0 8192 0 0 29 42 0 3
630 811
630 846
726 846
0 1 23 0 0 4096 0 0 44 38 0 3
700 828
700 877
731 877
0 1 23 0 0 12288 0 0 29 39 0 4
626 793
656 793
656 828
726 828
0 1 23 0 0 0 0 0 34 46 0 3
626 760
626 793
660 793
2 0 18 0 0 8320 0 32 0 0 134 3
668 1095
521 1095
521 552
2 0 20 0 0 8320 0 33 0 0 135 3
662 958
514 958
514 546
2 0 22 0 0 8320 0 34 0 0 136 3
660 811
509 811
509 523
1 0 17 0 0 8320 0 23 0 0 137 3
679 1192
462 1192
462 401
0 1 19 0 0 4224 0 0 24 138 0 3
476 287
476 1046
668 1046
0 1 21 0 0 4224 0 0 26 139 0 3
486 280
486 905
664 905
1 0 23 0 0 8320 0 25 0 0 140 3
660 760
500 760
500 236
5 2 24 0 0 8320 0 46 25 0 0 4
815 859
791 859
791 760
696 760
3 6 25 0 0 4224 0 34 46 0 0 4
709 802
807 802
807 868
815 868
7 3 26 0 0 8320 0 46 29 0 0 4
815 877
781 877
781 837
771 837
5 2 27 0 0 4224 0 42 26 0 0 4
819 999
716 999
716 905
700 905
3 6 28 0 0 4224 0 33 42 0 0 4
711 949
811 949
811 1008
819 1008
7 3 29 0 0 8320 0 42 30 0 0 4
819 1017
789 1017
789 978
779 978
2 5 30 0 0 4224 0 24 40 0 0 4
704 1046
802 1046
802 1139
820 1139
3 6 31 0 0 4224 0 32 40 0 0 4
717 1086
807 1086
807 1148
820 1148
3 7 32 0 0 8320 0 28 40 0 0 4
789 1118
812 1118
812 1157
820 1157
5 2 33 0 0 8320 0 38 23 0 0 4
824 1290
739 1290
739 1192
715 1192
6 3 34 0 0 4224 0 38 31 0 0 4
824 1299
733 1299
733 1232
725 1232
7 3 35 0 0 8320 0 38 27 0 0 4
824 1308
803 1308
803 1270
801 1270
8 3 36 0 0 4224 0 38 35 0 0 4
824 1317
800 1317
800 1320
799 1320
8 3 37 0 0 4224 0 40 36 0 0 2
820 1166
793 1166
8 3 38 0 0 4224 0 42 37 0 0 2
819 1026
785 1026
3 8 39 0 0 4224 0 44 46 0 0 2
777 886
815 886
12 0 40 0 0 4096 0 38 0 0 91 4
888 1281
929 1281
929 1282
934 1282
11 0 41 0 0 4096 0 38 0 0 92 2
888 1272
914 1272
12 0 40 0 0 4096 0 40 0 0 91 2
884 1130
934 1130
11 0 41 0 0 4096 0 40 0 0 92 2
884 1121
914 1121
12 0 40 0 0 4096 0 42 0 0 91 2
883 990
934 990
11 0 41 0 0 4096 0 42 0 0 92 2
883 981
914 981
10 0 2 0 0 4096 0 38 0 0 70 4
888 1263
905 1263
905 1254
908 1254
9 1 2 0 0 4096 0 38 39 0 0 3
894 1254
954 1254
954 1258
10 0 2 0 0 0 0 40 0 0 72 4
884 1112
901 1112
901 1103
904 1103
9 1 2 0 0 4096 0 40 41 0 0 3
890 1103
952 1103
952 1106
10 0 2 0 0 0 0 42 0 0 74 4
883 972
898 972
898 963
901 963
9 1 2 0 0 0 0 42 43 0 0 3
889 963
949 963
949 967
0 9 2 0 0 0 0 0 46 76 0 3
886 832
886 823
885 823
10 1 2 0 0 0 0 46 45 0 0 4
879 832
886 832
886 833
945 833
11 0 41 0 0 0 0 46 0 0 92 4
879 841
908 841
908 842
913 842
12 0 40 0 0 4096 0 46 0 0 91 2
879 850
934 850
8 13 42 0 0 4224 0 72 52 0 0 4
1001 707
886 707
886 696
872 696
0 1 7 0 0 0 0 0 47 126 0 2
1135 689
1135 676
4 1 23 0 0 0 0 69 12 0 0 6
1001 231
910 231
910 178
572 178
572 214
563 214
3 0 8 0 0 0 0 62 0 0 83 3
1175 508
1175 519
1125 519
10 1 8 0 0 0 0 71 66 0 0 3
1064 519
1125 519
1125 509
1 10 9 0 0 0 0 67 70 0 0 3
1123 364
1123 378
1066 378
11 0 41 0 0 4096 0 52 0 0 92 2
872 660
911 660
12 0 40 0 0 4096 0 52 0 0 91 2
872 669
934 669
12 0 40 0 0 4096 0 53 0 0 91 2
868 528
934 528
11 0 41 0 0 0 0 54 0 0 92 4
864 393
881 393
881 392
911 392
11 0 41 0 0 4096 0 53 0 0 92 2
868 519
911 519
12 0 40 0 0 4096 0 54 0 0 91 2
864 402
934 402
1 12 40 0 0 8320 0 2 55 0 0 5
962 1360
934 1360
934 260
862 260
862 248
1 11 41 0 0 12416 0 3 55 0 0 11
914 1359
914 1361
914 1361
914 842
913 842
913 660
911 660
911 249
866 249
866 239
862 239
8 13 43 0 0 4224 0 71 53 0 0 4
1000 537
874 537
874 555
868 555
8 13 44 0 0 4224 0 70 54 0 0 4
1002 396
878 396
878 429
864 429
13 8 45 0 0 4224 0 55 69 0 0 4
862 275
949 275
949 267
1001 267
10 0 2 0 0 0 0 52 0 0 97 3
872 651
881 651
881 641
9 1 2 0 0 12288 0 52 48 0 0 5
878 642
881 642
881 641
945 641
945 647
10 0 2 0 0 0 0 53 0 0 99 3
868 510
880 510
880 501
9 1 2 0 0 0 0 53 49 0 0 3
874 501
898 501
898 504
10 0 2 0 0 0 0 54 0 0 101 3
864 384
881 384
881 375
1 9 2 0 0 0 0 50 54 0 0 3
894 379
894 375
870 375
9 0 2 0 0 0 0 55 0 0 103 3
868 221
868 221
884 222
10 1 2 0 0 0 0 55 51 0 0 5
862 230
884 230
884 222
897 222
897 230
5 0 46 0 0 4096 0 52 0 0 124 4
808 678
780 678
780 677
765 677
7 0 16 0 0 0 0 52 0 0 123 3
808 696
664 696
664 669
0 7 18 0 0 0 0 0 53 120 0 3
656 518
656 555
804 555
0 7 20 0 0 0 0 0 54 135 0 2
671 429
800 429
0 7 22 0 0 0 0 0 55 122 0 3
660 244
660 275
798 275
6 2 47 0 0 4224 0 55 59 0 0 4
798 266
718 266
718 244
705 244
6 2 48 0 0 4224 0 54 58 0 0 4
800 420
718 420
718 406
710 406
2 6 49 0 0 4224 0 57 53 0 0 4
716 518
788 518
788 546
804 546
2 6 50 0 0 4224 0 56 52 0 0 4
712 669
791 669
791 687
808 687
5 0 46 0 0 4096 0 53 0 0 124 2
804 537
728 537
5 0 46 0 0 0 0 54 0 0 124 2
800 411
728 411
5 0 46 0 0 0 0 55 0 0 124 2
798 257
728 257
8 0 2 0 0 0 0 53 0 0 119 4
804 564
756 564
756 565
751 565
8 0 2 0 0 0 0 54 0 0 119 2
800 438
751 438
0 8 2 0 0 0 0 0 55 119 0 2
751 284
798 284
1 8 2 0 0 12416 0 60 52 0 0 5
769 128
769 130
751 130
751 705
808 705
1 0 18 0 0 0 0 57 0 0 134 4
680 518
574 518
574 554
575 554
0 1 20 0 0 0 0 0 7 135 0 2
567 536
566 536
1 1 22 0 0 0 0 8 59 0 0 4
563 480
598 480
598 244
669 244
0 1 16 0 0 0 0 0 56 133 0 2
584 669
676 669
2 0 46 0 0 4224 0 61 0 0 0 3
728 131
728 677
772 677
1 11 51 0 0 12416 0 63 72 0 0 5
1137 747
1137 759
1080 759
1080 680
1065 680
10 4 7 0 0 0 0 72 62 0 0 3
1065 689
1169 689
1169 508
0 2 9 0 0 0 0 0 62 84 0 7
1123 378
1134 378
1134 377
1150 377
1150 513
1181 513
1181 508
0 1 10 0 0 0 0 0 62 130 0 5
1121 247
1121 328
1200 328
1200 508
1187 508
11 9 52 0 0 8320 0 71 72 0 0 5
1064 510
1097 510
1097 748
1001 748
1001 716
10 1 10 0 0 0 0 69 68 0 0 3
1065 249
1121 249
1121 196
11 9 53 0 0 8320 0 70 71 0 0 5
1066 369
1082 369
1082 564
1000 564
1000 546
11 9 54 0 0 8320 0 69 70 0 0 5
1065 240
1075 240
1075 418
1002 418
1002 405
1 4 16 0 0 0 0 5 64 0 0 5
562 669
584 669
584 561
419 561
419 508
1 3 18 0 0 0 0 6 64 0 0 5
565 597
575 597
575 552
425 552
425 508
1 2 20 0 0 0 0 58 64 0 0 7
674 406
671 406
671 536
567 536
567 546
431 546
431 508
1 1 22 0 0 0 0 8 64 0 0 5
563 480
564 480
564 523
437 523
437 508
1 4 17 0 0 0 0 9 65 0 0 5
565 401
437 401
437 298
438 298
438 227
0 3 19 0 0 0 0 0 65 142 0 4
582 342
582 287
444 287
444 227
0 2 21 0 0 0 0 0 65 143 0 3
564 280
450 280
450 227
1 1 23 0 0 0 0 12 65 0 0 5
563 214
572 214
572 236
456 236
456 227
1 4 17 0 0 0 0 9 72 0 0 5
565 401
565 465
970 465
970 671
1001 671
1 4 19 0 0 0 0 10 71 0 0 4
563 342
963 342
963 501
1000 501
1 4 21 0 0 0 0 11 70 0 0 5
564 269
564 319
968 319
968 360
1002 360
1 9 55 0 0 4224 0 4 69 0 0 4
561 154
969 154
969 276
1001 276
35
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1288 926 1336 949
1301 936 1322 951
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1238 910 1349 933
1251 920 1335 935
12 Final Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
957 810 1066 833
969 820 1053 835
12 Logic Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1060 122 1204 145
1072 132 1191 147
17 Arithmetic Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
996 829 1044 852
1009 839 1030 854
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 32
691 1492 936 1515
701 1502 925 1517
32 ARITHMETIC LOGIC UNIT (METHOD I)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
871 1438 910 1461
883 1448 897 1463
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 15
786 728 916 751
798 738 903 753
15 ARITHMETIC UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 10
792 1364 887 1387
804 1374 874 1389
10 LOGIC UNIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
968 202 1007 225
980 212 994 227
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
897 1387 936 1410
909 1397 923 1412
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
951 1388 992 1411
964 1398 978 1413
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
428 421 463 444
441 431 449 446
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
424 128 459 151
437 138 445 153
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1138 170 1186 193
1151 180 1172 195
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
979 747 1090 770
992 757 1076 772
12 Full Adder 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
989 563 1100 586
1002 573 1086 588
12 Full Adder 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
986 413 1095 436
998 423 1082 438
12 Full Adder 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
976 278 1085 301
988 288 1072 303
12 Full Adder 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
976 676 1015 699
988 686 1002 701
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
973 507 1014 530
986 517 1000 532
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
972 365 1013 388
985 375 999 390
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
974 237 1013 260
986 247 1000 262
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
473 392 512 415
485 402 499 417
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 322 512 345
484 332 498 347
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 258 510 281
483 268 497 283
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
470 193 509 216
482 203 496 218
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
475 462 516 485
488 472 502 487
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
477 523 518 546
490 533 504 548
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 580 518 603
491 590 505 605
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 657 518 680
491 667 505 682
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
461 141 509 164
474 151 495 166
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
972 637 1013 660
985 647 999 662
2 X3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
973 469 1012 492
985 479 999 494
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
972 332 1013 355
985 342 999 357
2 X1
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
