CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
450 740 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
76
13 Logic Switch~
5 943 1520 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
363 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 549 157 0 1 11
0 63
0
0 0 21360 0
2 0V
-8 -17 6 -9
3 V11
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8132 0 0
2
43336.5 0
0
13 Logic Switch~
5 550 669 0 1 11
0 14
0
0 0 21360 0
2 0V
-8 -16 6 -8
3 V10
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
65 0 0
2
5.89859e-315 5.26354e-315
0
13 Logic Switch~
5 553 597 0 1 11
0 15
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
6609 0 0
2
5.89859e-315 5.30499e-315
0
13 Logic Switch~
5 552 536 0 1 11
0 16
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V8
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8995 0 0
2
5.89859e-315 5.32571e-315
0
13 Logic Switch~
5 551 480 0 1 11
0 17
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3918 0 0
2
5.89859e-315 5.34643e-315
0
13 Logic Switch~
5 553 401 0 1 11
0 18
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7519 0 0
2
5.89859e-315 5.3568e-315
0
13 Logic Switch~
5 551 342 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
377 0 0
2
5.89859e-315 5.36716e-315
0
13 Logic Switch~
5 552 269 0 1 11
0 19
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
8816 0 0
2
5.89859e-315 5.37752e-315
0
13 Logic Switch~
5 551 214 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -19 7 -11
2 V3
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3877 0 0
2
5.89859e-315 5.38788e-315
0
13 Logic Switch~
5 903 1447 0 1 11
0 38
0
0 0 21360 90
2 0V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
926 0 0
2
5.89859e-315 5.39306e-315
0
13 Logic Switch~
5 960 1444 0 1 11
0 39
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7262 0 0
2
5.89859e-315 5.39824e-315
0
14 Logic Display~
6 1016 1260 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L19
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5267 0 0
2
43336.5 0
0
7 Ground~
168 1133 1215 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8838 0 0
2
43336.5 0
0
14 Logic Display~
6 1316 1304 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7159 0 0
2
43336.5 0
0
7 74LS157
122 1167 1147 0 14 29
0 12 42 7 13 6 3 5 40 4
2 11 10 9 8
0
0 0 4848 0
7 74LS157
-24 -60 25 -52
2 U8
-7 -61 7 -53
0
15 DVCC=16;DGND=8;
131 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 2 6 5 10 11 13 14
15 4 7 9 12 1 3 2 6 5
10 11 13 14 15 4 7 9 12 0
65 0 0 0 0 0 0 0
1 U
5812 0 0
2
43336.5 0
0
5 4071~
219 761 1420 0 3 22
0 18 14 25
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U21C
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 9 0
1 U
331 0 0
2
5.89859e-315 5.40342e-315
0
5 4030~
219 687 1344 0 3 22
0 18 14 23
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U18D
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 6 0
1 U
9604 0 0
2
5.89859e-315 5.4086e-315
0
5 4081~
219 767 1363 0 3 22
0 18 14 24
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19D
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 7 0
1 U
7518 0 0
2
5.89859e-315 5.41378e-315
0
5 4069~
219 687 1299 0 2 22
0 18 22
0
0 0 624 0
4 4069
-7 -24 21 -16
4 U20D
-14 -20 14 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 8 0
1 U
4832 0 0
2
5.89859e-315 5.41896e-315
0
5 4071~
219 757 1264 0 3 22
0 20 15 29
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U21B
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 9 0
1 U
6798 0 0
2
5.89859e-315 5.42414e-315
0
5 4030~
219 683 1188 0 3 22
0 20 15 27
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U18C
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 6 0
1 U
3336 0 0
2
5.89859e-315 5.42933e-315
0
5 4081~
219 763 1207 0 3 22
0 20 15 28
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 7 0
1 U
8370 0 0
2
5.89859e-315 5.43192e-315
0
5 4069~
219 683 1143 0 2 22
0 20 26
0
0 0 624 0
4 4069
-7 -24 21 -16
4 U20C
-14 -20 14 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 8 0
1 U
3910 0 0
2
5.89859e-315 5.43451e-315
0
5 4071~
219 755 1105 0 3 22
0 19 16 33
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U21A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 9 0
1 U
316 0 0
2
5.89859e-315 5.4371e-315
0
5 4030~
219 681 1029 0 3 22
0 19 16 31
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U18B
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 6 0
1 U
536 0 0
2
5.89859e-315 5.43969e-315
0
5 4081~
219 761 1048 0 3 22
0 19 16 32
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 7 0
1 U
4460 0 0
2
5.89859e-315 5.44228e-315
0
5 4069~
219 681 984 0 2 22
0 19 30
0
0 0 624 0
4 4069
-7 -24 21 -16
4 U20B
-14 -20 14 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 8 0
1 U
3260 0 0
2
5.89859e-315 5.44487e-315
0
5 4069~
219 676 821 0 2 22
0 21 34
0
0 0 624 0
4 4069
-7 -24 21 -16
4 U20A
-14 -20 14 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 8 0
1 U
5156 0 0
2
5.89859e-315 5.44746e-315
0
5 4081~
219 756 885 0 3 22
0 21 17 36
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U19A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 7 0
1 U
3133 0 0
2
5.89859e-315 5.45005e-315
0
5 4030~
219 676 866 0 3 22
0 21 17 35
0
0 0 624 0
4 4030
-7 -24 21 -16
4 U18A
-8 -25 20 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
5523 0 0
2
5.89859e-315 5.45264e-315
0
5 4071~
219 750 942 0 3 22
0 21 17 37
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U17A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3746 0 0
2
5.89859e-315 5.45523e-315
0
7 74LS151
20 847 1362 0 14 29
0 64 65 66 67 22 23 24 25 2
2 38 39 40 68
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U16
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
5668 0 0
2
5.89859e-315 5.45782e-315
0
7 Ground~
168 906 1345 0 1 3
0 2
0
0 0 53360 0
0
4 GND9
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
5368 0 0
2
5.89859e-315 5.46041e-315
0
7 Ground~
168 903 1188 0 1 3
0 2
0
0 0 53360 0
0
4 GND7
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
8293 0 0
2
5.89859e-315 5.463e-315
0
7 74LS151
20 844 1205 0 14 29
0 69 70 71 72 26 27 28 29 2
2 38 39 3 73
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U15
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
3232 0 0
2
5.89859e-315 5.46559e-315
0
14 Logic Display~
6 1015 1327 0 1 2
10 41
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L15
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6644 0 0
2
5.89859e-315 5.46818e-315
0
14 Logic Display~
6 1001 1036 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L13
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4978 0 0
2
5.89859e-315 5.47207e-315
0
7 74LS151
20 841 1047 0 14 29
0 74 75 76 77 30 31 32 33 2
2 38 39 13 78
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U14
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
9207 0 0
2
5.89859e-315 5.47336e-315
0
7 Ground~
168 899 1032 0 1 3
0 2
0
0 0 53360 0
0
4 GND6
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
6998 0 0
2
5.89859e-315 5.47466e-315
0
14 Logic Display~
6 998 865 0 1 2
10 42
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L12
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3175 0 0
2
5.89859e-315 5.47595e-315
0
7 Ground~
168 896 869 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3378 0 0
2
5.89859e-315 5.47725e-315
0
7 74LS151
20 838 884 0 14 29
0 79 80 81 82 34 35 36 37 2
2 38 39 42 83
0
0 0 4848 0
7 74LS151
-24 -60 25 -52
3 U13
-10 -61 11 -53
0
15 DVCC=16;DGND=8;
141 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i %10i %11i %12i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 12 13 14 15 1 2 3 4 7
9 10 11 5 6 12 13 14 15 1
2 3 4 7 9 10 11 5 6 0
65 0 0 512 1 0 0 0
1 U
922 0 0
2
5.89859e-315 5.47854e-315
0
14 Logic Display~
6 1314 1233 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6891 0 0
2
5.89859e-315 5.48113e-315
0
14 Logic Display~
6 1311 1166 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5407 0 0
2
5.89859e-315 5.48502e-315
0
14 Logic Display~
6 1308 1110 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7349 0 0
2
5.89859e-315 5.4889e-315
0
5 4049~
219 816 748 0 2 22
0 14 43
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
3919 0 0
2
43336.5 1
0
5 4049~
219 818 586 0 2 22
0 15 44
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
9747 0 0
2
43336.5 2
0
12 Hex Display~
7 1420 476 0 18 19
10 7 6 5 4 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
5310 0 0
2
43336.5 3
0
14 Logic Display~
6 1295 780 0 1 2
10 47
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4318 0 0
2
43336.5 4
0
12 Hex Display~
7 400 491 0 16 19
10 17 16 15 14 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3917 0 0
2
43336.5 5
0
12 Hex Display~
7 396 207 0 18 19
10 21 19 20 18 0 0 0 0 0
0 1 0 1 1 0 1 1 5
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7930 0 0
2
43336.5 6
0
14 Logic Display~
6 1292 643 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6128 0 0
2
43336.5 7
0
14 Logic Display~
6 1292 483 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7346 0 0
2
43336.5 8
0
14 Logic Display~
6 1288 343 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8577 0 0
2
43336.5 9
0
14 Logic Display~
6 1284 187 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3372 0 0
2
43336.5 10
0
14 Logic Display~
6 731 130 0 1 2
10 39
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3741 0 0
2
43336.5 11
0
14 Logic Display~
6 685 131 0 1 2
10 38
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5813 0 0
2
43336.5 12
0
5 4071~
219 979 712 0 3 22
0 56 55 53
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
3213 0 0
2
43336.5 13
0
5 4071~
219 974 547 0 3 22
0 58 57 51
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
3694 0 0
2
43336.5 14
0
5 4071~
219 969 397 0 3 22
0 60 59 54
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4327 0 0
2
43336.5 15
0
5 4071~
219 962 242 0 3 22
0 61 62 52
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
8800 0 0
2
43336.5 16
0
5 4049~
219 806 432 0 2 22
0 16 46
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
3406 0 0
2
43336.5 17
0
5 4049~
219 800 285 0 2 22
0 17 45
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
6455 0 0
2
43336.5 18
0
4 4008
219 1148 216 0 14 29
0 84 85 86 21 87 88 89 52 63
7 50 90 91 92
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9319 0 0
2
5.89859e-315 5.49538e-315
0
4 4008
219 1154 370 0 14 29
0 93 94 95 19 96 97 98 54 50
6 49 99 100 101
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3172 0 0
2
5.89859e-315 5.49667e-315
0
4 4008
219 1151 521 0 14 29
0 102 103 104 20 105 106 107 51 49
5 48 108 109 110
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
38 0 0
2
5.89859e-315 5.49797e-315
0
4 4008
219 1152 686 0 14 29
0 111 112 113 18 114 115 116 53 48
4 47 117 118 119
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
376 0 0
2
5.89859e-315 5.49926e-315
0
5 4081~
219 866 210 0 3 22
0 39 17 61
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
6666 0 0
2
5.89859e-315 5.50056e-315
0
5 4081~
219 864 294 0 3 22
0 45 38 62
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
9365 0 0
2
5.89859e-315 5.50185e-315
0
5 4081~
219 866 367 0 3 22
0 39 16 60
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3251 0 0
2
5.89859e-315 5.50315e-315
0
5 4081~
219 868 441 0 3 22
0 46 38 59
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
5481 0 0
2
5.89859e-315 5.50444e-315
0
5 4081~
219 873 520 0 3 22
0 39 15 58
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
7788 0 0
2
5.89859e-315 5.50574e-315
0
5 4081~
219 875 595 0 3 22
0 44 38 57
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3273 0 0
2
5.89859e-315 5.50703e-315
0
5 4081~
219 874 683 0 3 22
0 39 14 56
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3761 0 0
2
5.89859e-315 5.50833e-315
0
5 4081~
219 872 757 0 3 22
0 43 38 55
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3226 0 0
2
5.89859e-315 5.50963e-315
0
139
1 0 3 0 0 12288 0 13 0 0 66 4
1016 1278
1016 1282
978 1282
978 1232
0 9 4 0 0 4224 0 0 16 98 0 5
1345 694
1345 1044
1094 1044
1094 1183
1135 1183
0 7 5 0 0 4224 0 0 16 99 0 5
1366 527
1366 1064
1078 1064
1078 1165
1135 1165
0 5 6 0 0 4224 0 0 16 100 0 5
1394 513
1394 1086
1101 1086
1101 1147
1135 1147
0 3 7 0 0 4224 0 0 16 101 0 5
1440 508
1440 1091
1106 1091
1106 1129
1135 1129
10 1 2 0 0 8192 0 16 14 0 0 5
1129 1192
1125 1192
1125 1201
1133 1201
1133 1209
1 14 8 0 0 12416 0 15 16 0 0 5
1316 1322
1316 1326
1207 1326
1207 1183
1199 1183
13 1 9 0 0 4224 0 16 44 0 0 5
1199 1165
1294 1165
1294 1259
1314 1259
1314 1251
12 1 10 0 0 4224 0 16 45 0 0 5
1199 1147
1298 1147
1298 1192
1311 1192
1311 1184
11 1 11 0 0 4224 0 16 46 0 0 3
1199 1129
1308 1129
1308 1128
1 1 12 0 0 8320 0 1 16 0 0 4
955 1520
1121 1520
1121 1111
1135 1111
13 4 13 0 0 4224 0 39 16 0 0 5
873 1074
1111 1074
1111 1139
1135 1139
1135 1138
0 2 14 0 0 4096 0 0 17 14 0 3
709 1372
709 1429
748 1429
0 2 14 0 0 8192 0 0 19 21 0 3
661 1353
661 1372
743 1372
0 2 15 0 0 4096 0 0 21 16 0 3
709 1216
709 1273
744 1273
0 2 15 0 0 8192 0 0 23 22 0 3
655 1197
655 1216
739 1216
0 2 16 0 0 4096 0 0 25 18 0 3
724 1057
724 1114
742 1114
0 2 16 0 0 8192 0 0 27 23 0 3
657 1038
657 1057
737 1057
0 2 17 0 0 4096 0 0 32 20 0 3
682 894
682 951
737 951
0 2 17 0 0 8192 0 0 30 24 0 3
620 875
620 894
732 894
2 0 14 0 0 8320 0 18 0 0 87 3
671 1353
573 1353
573 722
2 0 15 0 0 8320 0 22 0 0 110 3
667 1197
419 1197
419 552
2 0 16 0 0 8320 0 26 0 0 111 3
665 1038
427 1038
427 546
0 2 17 0 0 4224 0 0 31 112 0 3
437 523
437 875
660 875
1 0 18 0 0 8192 0 17 0 0 26 3
748 1411
724 1411
724 1364
0 1 18 0 0 8192 0 0 19 27 0 5
645 1335
645 1364
735 1364
735 1354
743 1354
1 0 18 0 0 0 0 18 0 0 37 3
671 1335
645 1335
645 1299
1 0 19 0 0 8192 0 25 0 0 29 3
742 1096
706 1096
706 1049
0 1 19 0 0 8192 0 0 27 33 0 5
647 1020
647 1049
729 1049
729 1039
737 1039
0 1 20 0 0 4096 0 0 21 31 0 3
727 1208
727 1255
744 1255
0 1 20 0 0 12288 0 0 23 32 0 6
641 1177
642 1177
642 1208
731 1208
731 1198
739 1198
0 1 20 0 0 0 0 0 22 38 0 3
641 1143
641 1179
667 1179
0 1 19 0 0 0 0 0 26 39 0 3
647 984
647 1020
665 1020
0 1 21 0 0 4096 0 0 32 35 0 3
710 886
710 933
737 933
0 1 21 0 0 8192 0 0 30 36 0 5
637 857
637 886
724 886
724 876
732 876
0 1 21 0 0 0 0 0 31 40 0 3
634 821
634 857
660 857
0 1 18 0 0 4224 0 0 20 113 0 3
456 401
456 1299
672 1299
1 0 20 0 0 8320 0 24 0 0 114 3
668 1143
473 1143
473 287
0 1 19 0 0 4224 0 0 28 115 0 3
491 280
491 984
666 984
0 1 21 0 0 4224 0 0 29 116 0 3
504 242
504 821
661 821
2 5 22 0 0 4224 0 20 33 0 0 4
708 1299
799 1299
799 1371
815 1371
3 6 23 0 0 4224 0 18 33 0 0 4
720 1344
804 1344
804 1380
815 1380
3 7 24 0 0 8320 0 19 33 0 0 4
788 1363
809 1363
809 1389
815 1389
3 8 25 0 0 8320 0 17 33 0 0 4
794 1420
809 1420
809 1398
815 1398
2 5 26 0 0 4224 0 24 36 0 0 5
704 1143
795 1143
795 1215
812 1215
812 1214
3 6 27 0 0 4224 0 22 36 0 0 5
716 1188
800 1188
800 1224
812 1224
812 1223
3 7 28 0 0 8320 0 23 36 0 0 5
784 1207
805 1207
805 1233
812 1233
812 1232
3 8 29 0 0 8320 0 21 36 0 0 5
790 1264
805 1264
805 1242
812 1242
812 1241
2 5 30 0 0 4224 0 28 39 0 0 4
702 984
793 984
793 1056
809 1056
3 6 31 0 0 4224 0 26 39 0 0 4
714 1029
798 1029
798 1065
809 1065
3 7 32 0 0 8320 0 27 39 0 0 4
782 1048
803 1048
803 1074
809 1074
3 8 33 0 0 8320 0 25 39 0 0 4
788 1105
803 1105
803 1083
809 1083
2 5 34 0 0 4224 0 29 43 0 0 4
697 821
788 821
788 893
806 893
3 6 35 0 0 4224 0 31 43 0 0 4
709 866
793 866
793 902
806 902
3 7 36 0 0 8320 0 30 43 0 0 4
777 885
798 885
798 911
806 911
3 8 37 0 0 8320 0 32 43 0 0 4
783 942
798 942
798 920
806 920
11 0 38 0 0 4096 0 43 0 0 139 2
870 875
928 875
12 0 39 0 0 4096 0 43 0 0 138 2
870 884
968 884
11 0 38 0 0 0 0 39 0 0 139 2
873 1038
928 1038
12 0 39 0 0 0 0 39 0 0 138 2
873 1047
968 1047
11 0 38 0 0 0 0 36 0 0 139 4
876 1196
890 1196
890 1197
928 1197
12 0 39 0 0 0 0 36 0 0 138 2
876 1205
968 1205
0 11 38 0 0 0 0 0 33 139 0 4
928 1354
893 1354
893 1353
879 1353
12 0 39 0 0 0 0 33 0 0 138 2
879 1362
968 1362
8 13 40 0 0 12416 0 16 33 0 0 4
1135 1174
1109 1174
1109 1389
879 1389
6 13 3 0 0 12416 0 16 36 0 0 4
1135 1156
1114 1156
1114 1232
876 1232
0 1 41 0 0 4224 0 0 37 0 0 2
1015 1389
1015 1345
10 0 2 0 0 4096 0 33 0 0 69 3
879 1344
892 1344
892 1335
1 9 2 0 0 12416 0 34 33 0 0 4
906 1339
905 1339
905 1335
885 1335
10 0 2 0 0 0 0 36 0 0 71 3
876 1187
889 1187
889 1178
1 9 2 0 0 0 0 35 36 0 0 4
903 1182
902 1182
902 1178
882 1178
1 0 13 0 0 128 0 38 0 0 12 2
1001 1054
1001 1074
10 0 2 0 0 0 0 39 0 0 74 3
873 1029
886 1029
886 1020
1 9 2 0 0 0 0 40 39 0 0 3
899 1026
899 1020
879 1020
0 1 42 0 0 4096 0 0 41 76 0 2
998 911
998 883
13 2 42 0 0 4224 0 43 16 0 0 4
870 911
1116 911
1116 1120
1135 1120
10 0 2 0 0 0 0 43 0 0 78 3
870 866
883 866
883 857
1 9 2 0 0 0 0 42 43 0 0 3
896 863
896 857
876 857
2 0 38 0 0 4096 0 76 0 0 139 2
848 766
683 766
1 0 39 0 0 4096 0 75 0 0 138 2
850 674
730 674
0 0 38 0 0 0 0 0 0 136 139 2
834 604
683 604
1 0 39 0 0 0 0 73 0 0 138 2
849 511
730 511
2 0 38 0 0 0 0 72 0 0 139 2
844 450
683 450
1 0 39 0 0 0 0 71 0 0 138 4
842 358
736 358
736 359
730 359
2 0 38 0 0 0 0 70 0 0 139 2
840 303
683 303
1 0 39 0 0 0 0 69 0 0 138 2
842 201
730 201
0 1 14 0 0 0 0 0 3 89 0 4
786 722
573 722
573 669
562 669
1 0 14 0 0 0 0 47 0 0 89 4
801 748
793 748
793 747
786 747
2 0 14 0 0 0 0 75 0 0 0 4
850 692
786 692
786 747
781 747
1 2 43 0 0 4224 0 76 47 0 0 2
848 748
837 748
0 2 15 0 0 0 0 0 73 123 0 4
786 560
785 560
785 529
849 529
1 2 44 0 0 4224 0 74 48 0 0 2
851 586
839 586
2 0 16 0 0 0 0 71 0 0 124 3
842 376
783 376
783 399
0 2 17 0 0 0 0 0 69 125 0 3
777 249
777 219
842 219
1 2 45 0 0 4224 0 70 64 0 0 2
840 285
821 285
1 2 46 0 0 4224 0 72 63 0 0 2
844 432
827 432
1 11 47 0 0 12416 0 50 68 0 0 5
1295 798
1295 802
1192 802
1192 686
1184 686
0 4 4 0 0 0 0 0 49 102 0 3
1292 694
1411 694
1411 500
0 3 5 0 0 0 0 0 49 104 0 3
1292 527
1417 527
1417 500
0 2 6 0 0 0 0 0 49 105 0 6
1288 379
1288 444
1375 444
1375 513
1423 513
1423 500
0 1 7 0 0 0 0 0 49 106 0 6
1284 225
1284 328
1449 328
1449 508
1429 508
1429 500
1 10 4 0 0 0 0 53 68 0 0 3
1292 661
1292 695
1184 695
11 9 48 0 0 8320 0 67 68 0 0 6
1183 521
1188 521
1188 737
1112 737
1112 722
1120 722
1 10 5 0 0 0 0 54 67 0 0 3
1292 501
1292 530
1183 530
10 1 6 0 0 0 0 66 55 0 0 3
1186 379
1288 379
1288 361
10 1 7 0 0 0 0 65 56 0 0 3
1180 225
1284 225
1284 205
11 9 49 0 0 8320 0 66 67 0 0 6
1186 370
1195 370
1195 572
1111 572
1111 557
1119 557
11 9 50 0 0 8320 0 65 66 0 0 6
1180 216
1190 216
1190 421
1114 421
1114 406
1122 406
0 4 14 0 0 0 0 0 51 87 0 5
573 669
575 669
575 558
391 558
391 515
1 3 15 0 0 0 0 4 51 0 0 5
565 597
575 597
575 552
397 552
397 515
0 2 16 0 0 0 0 0 51 124 0 4
567 536
567 546
403 546
403 515
0 1 17 0 0 0 0 0 51 125 0 4
569 480
569 523
409 523
409 515
1 4 18 0 0 0 0 7 52 0 0 5
565 401
388 401
388 298
387 298
387 231
0 3 20 0 0 0 0 0 52 118 0 4
582 342
582 287
393 287
393 231
0 2 19 0 0 0 0 0 52 119 0 3
564 280
399 280
399 231
1 1 21 0 0 0 0 10 52 0 0 5
563 214
564 214
564 242
405 242
405 231
1 4 18 0 0 0 0 7 68 0 0 5
565 401
565 465
1015 465
1015 677
1120 677
1 4 20 0 0 0 0 8 67 0 0 4
563 342
1110 342
1110 512
1119 512
1 4 19 0 0 0 0 9 66 0 0 5
564 269
564 319
1092 319
1092 361
1122 361
1 4 21 0 0 0 0 10 65 0 0 6
563 214
564 214
564 181
1075 181
1075 207
1116 207
3 8 51 0 0 4224 0 60 67 0 0 4
1007 547
1110 547
1110 548
1119 548
3 8 52 0 0 4224 0 62 65 0 0 4
995 242
1080 242
1080 243
1116 243
1 1 15 0 0 0 0 4 48 0 0 6
565 597
589 597
589 560
786 560
786 586
803 586
1 1 16 0 0 0 0 5 63 0 0 6
564 536
591 536
591 399
783 399
783 432
791 432
1 1 17 0 0 0 0 6 64 0 0 6
563 480
617 480
617 249
778 249
778 285
785 285
3 8 53 0 0 4224 0 59 68 0 0 4
1012 712
1096 712
1096 713
1120 713
3 8 54 0 0 4224 0 61 66 0 0 2
1002 397
1122 397
2 3 55 0 0 4224 0 59 76 0 0 4
966 721
901 721
901 757
893 757
1 3 56 0 0 4224 0 59 75 0 0 4
966 703
903 703
903 683
895 683
2 3 57 0 0 4224 0 60 74 0 0 4
961 556
904 556
904 595
896 595
1 3 58 0 0 4224 0 60 73 0 0 4
961 538
902 538
902 520
894 520
2 3 59 0 0 4224 0 61 72 0 0 4
956 406
897 406
897 441
889 441
1 3 60 0 0 4224 0 61 71 0 0 4
956 388
895 388
895 367
887 367
3 1 61 0 0 4224 0 69 62 0 0 4
887 210
940 210
940 233
949 233
3 2 62 0 0 4224 0 70 62 0 0 4
885 294
940 294
940 251
949 251
2 0 38 0 0 0 0 74 0 0 0 2
851 604
830 604
1 9 63 0 0 4224 0 2 65 0 0 4
561 157
1070 157
1070 252
1116 252
1 1 39 0 0 24704 0 12 57 0 0 8
961 1431
967 1431
967 1407
968 1407
968 796
730 796
730 148
731 148
1 1 38 0 0 12416 0 11 58 0 0 7
904 1434
904 1427
928 1427
928 781
683 781
683 149
685 149
35
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
384 418 419 441
397 428 405 443
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
379 131 414 154
392 141 400 156
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1296 199 1344 222
1309 209 1330 224
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1098 742 1209 765
1111 752 1195 767
12 Full Adder 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1096 570 1207 593
1109 580 1193 595
12 Full Adder 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1100 421 1209 444
1112 431 1196 446
12 Full Adder 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1096 264 1205 287
1108 274 1192 289
12 Full Adder 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1081 710 1120 733
1093 720 1107 735
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1077 545 1118 568
1090 555 1104 570
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1076 394 1117 417
1089 404 1103 419
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1085 216 1124 239
1097 226 1111 241
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
473 392 512 415
485 402 499 417
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 322 512 345
484 332 498 347
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 258 510 281
483 268 497 283
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
470 193 509 216
482 203 496 218
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
475 462 516 485
488 472 502 487
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
477 523 518 546
490 533 504 548
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 580 518 603
491 590 505 605
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 657 518 680
491 667 505 682
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
461 141 509 164
474 151 495 166
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1083 649 1124 672
1096 659 1110 674
2 X3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1076 499 1115 522
1088 509 1102 524
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1077 357 1118 380
1090 367 1104 382
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1084 189 1123 212
1096 199 1110 214
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
944 1452 985 1475
957 1462 971 1477
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
880 1459 919 1482
892 1469 906 1484
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
919 1529 960 1552
932 1539 946 1554
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 18
1007 776 1158 799
1019 786 1145 801
18 ARITHMETIC CIRCUIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 13
783 1433 901 1456
796 1443 887 1458
13 LOGIC CIRCUIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 33
813 1572 1069 1595
825 1582 1056 1597
33 ARITHMETIC LOGIC UNIT (METHOD II)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1334 1109 1382 1132
1347 1119 1368 1134
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1014 862 1062 885
1027 872 1048 887
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1234 112 1380 135
1247 122 1366 137
17 Arithmetic Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
971 809 1080 832
983 819 1067 834
12 Logic Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1319 1095 1430 1118
1332 1105 1416 1120
12 Final Output
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
