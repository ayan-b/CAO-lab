CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
310 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
43
13 Logic Switch~
5 672 793 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3273 0 0
2
43336 0
0
13 Logic Switch~
5 716 796 0 1 11
0 2
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
3761 0 0
2
43336 0
0
13 Logic Switch~
5 549 157 0 1 11
0 36
0
0 0 21360 0
2 0V
-8 -17 6 -9
3 V11
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3226 0 0
2
43336 0
0
13 Logic Switch~
5 550 669 0 10 11
0 4 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
3 V10
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4244 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 553 597 0 1 11
0 6
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5225 0 0
2
5.89859e-315 5.26354e-315
0
13 Logic Switch~
5 552 536 0 1 11
0 8
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V8
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
768 0 0
2
5.89859e-315 5.30499e-315
0
13 Logic Switch~
5 551 480 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
5735 0 0
2
5.89859e-315 5.32571e-315
0
13 Logic Switch~
5 553 401 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5881 0 0
2
5.89859e-315 5.34643e-315
0
13 Logic Switch~
5 551 342 0 1 11
0 21
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3275 0 0
2
5.89859e-315 5.3568e-315
0
13 Logic Switch~
5 552 269 0 1 11
0 22
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4203 0 0
2
5.89859e-315 5.36716e-315
0
13 Logic Switch~
5 551 214 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-7 -19 7 -11
2 V3
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3440 0 0
2
5.89859e-315 5.37752e-315
0
13 Logic Switch~
5 903 1447 0 10 11
0 37 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
11 0 25 8
2 V1
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -1 0
1 V
9102 0 0
2
5.89859e-315 5.38788e-315
0
13 Logic Switch~
5 960 1444 0 1 11
0 38
0
0 0 21360 90
2 0V
11 0 25 8
2 V2
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 512 1 0 -2 0
1 V
5586 0 0
2
5.89859e-315 5.39306e-315
0
5 4049~
219 816 748 0 2 22
0 4 5
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
525 0 0
2
43336 1
0
5 4049~
219 818 586 0 2 22
0 6 7
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
6206 0 0
2
43336 2
0
12 Hex Display~
7 1357 474 0 18 19
10 16 15 14 13 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3418 0 0
2
43336 3
0
14 Logic Display~
6 1295 780 0 1 2
10 12
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9312 0 0
2
43336 4
0
12 Hex Display~
7 400 491 0 18 19
10 9 8 6 4 0 0 0 0 0
0 1 1 1 1 1 1 1 8
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7419 0 0
2
43336 5
0
12 Hex Display~
7 396 207 0 18 19
10 23 22 21 20 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
472 0 0
2
43336 6
0
14 Logic Display~
6 1292 643 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4714 0 0
2
43336 7
0
14 Logic Display~
6 1292 483 0 1 2
10 14
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9386 0 0
2
43336 8
0
14 Logic Display~
6 1288 343 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7610 0 0
2
43336 9
0
14 Logic Display~
6 1284 187 0 1 2
10 16
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3482 0 0
2
43336 10
0
14 Logic Display~
6 730 130 0 1 2
10 2
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3608 0 0
2
43336 11
0
14 Logic Display~
6 683 132 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6397 0 0
2
43336 12
0
5 4071~
219 979 712 0 3 22
0 29 28 26
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
3967 0 0
2
43336 13
0
5 4071~
219 974 547 0 3 22
0 31 30 24
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
8621 0 0
2
43336 14
0
5 4071~
219 969 397 0 3 22
0 33 32 27
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
8901 0 0
2
43336 15
0
5 4071~
219 962 242 0 3 22
0 34 35 25
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
7385 0 0
2
43336 16
0
5 4049~
219 806 432 0 2 22
0 8 11
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7B
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
6519 0 0
2
43336 17
0
5 4049~
219 800 285 0 2 22
0 9 10
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
552 0 0
2
43336 18
0
4 4008
219 1148 216 0 14 29
0 39 40 41 23 42 43 44 25 36
16 19 45 46 47
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
5551 0 0
2
5.89859e-315 5.39824e-315
0
4 4008
219 1154 370 0 14 29
0 48 49 50 22 51 52 53 27 19
15 18 54 55 56
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8715 0 0
2
5.89859e-315 5.40342e-315
0
4 4008
219 1151 521 0 14 29
0 57 58 59 21 60 61 62 24 18
14 17 63 64 65
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9763 0 0
2
5.89859e-315 5.4086e-315
0
4 4008
219 1152 686 0 14 29
0 66 67 68 20 69 70 71 26 17
13 12 72 73 74
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
8443 0 0
2
5.89859e-315 5.41378e-315
0
5 4081~
219 866 210 0 3 22
0 2 9 34
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
3719 0 0
2
5.89859e-315 5.41896e-315
0
5 4081~
219 864 294 0 3 22
0 10 3 35
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
8671 0 0
2
5.89859e-315 5.42414e-315
0
5 4081~
219 866 367 0 3 22
0 2 8 33
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
7168 0 0
2
5.89859e-315 5.42933e-315
0
5 4081~
219 868 441 0 3 22
0 11 3 32
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
49 0 0
2
5.89859e-315 5.43192e-315
0
5 4081~
219 873 520 0 3 22
0 2 6 31
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
6536 0 0
2
5.89859e-315 5.43451e-315
0
5 4081~
219 875 595 0 3 22
0 7 3 30
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3931 0 0
2
5.89859e-315 5.4371e-315
0
5 4081~
219 874 683 0 3 22
0 2 4 29
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
4390 0 0
2
5.89859e-315 5.43969e-315
0
5 4081~
219 872 757 0 3 22
0 5 3 28
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3242 0 0
2
5.89859e-315 5.44228e-315
0
61
1 1 2 0 0 8320 0 2 24 0 0 3
728 796
730 796
730 148
1 1 3 0 0 8320 0 1 25 0 0 3
684 793
683 793
683 150
2 0 3 0 0 0 0 43 0 0 2 2
848 766
683 766
1 0 2 0 0 0 0 42 0 0 1 2
850 674
730 674
0 0 3 0 0 0 0 0 0 60 2 2
834 604
683 604
1 0 2 0 0 0 0 40 0 0 1 2
849 511
730 511
2 0 3 0 0 0 0 39 0 0 2 2
844 450
683 450
1 0 2 0 0 0 0 38 0 0 1 4
842 358
736 358
736 359
730 359
2 0 3 0 0 0 0 37 0 0 2 2
840 303
683 303
1 0 2 0 0 0 0 36 0 0 1 2
842 201
730 201
0 1 4 0 0 4224 0 0 4 13 0 4
786 722
573 722
573 669
562 669
1 0 4 0 0 0 0 14 0 0 13 4
801 748
793 748
793 747
786 747
2 0 4 0 0 0 0 42 0 0 0 4
850 692
786 692
786 747
781 747
1 2 5 0 0 4224 0 43 14 0 0 2
848 748
837 748
0 2 6 0 0 12288 0 0 40 47 0 4
786 560
785 560
785 529
849 529
1 2 7 0 0 4224 0 41 15 0 0 2
851 586
839 586
2 0 8 0 0 4096 0 38 0 0 48 3
842 376
783 376
783 399
0 2 9 0 0 8192 0 0 36 49 0 3
777 249
777 219
842 219
1 2 10 0 0 4224 0 37 31 0 0 2
840 285
821 285
1 2 11 0 0 4224 0 39 30 0 0 2
844 432
827 432
1 11 12 0 0 12416 0 17 35 0 0 5
1295 798
1295 802
1192 802
1192 686
1184 686
0 4 13 0 0 8320 0 0 16 26 0 3
1292 694
1348 694
1348 498
0 3 14 0 0 4096 0 0 16 28 0 3
1292 527
1354 527
1354 498
0 2 15 0 0 12288 0 0 16 29 0 6
1288 379
1288 444
1322 444
1322 513
1360 513
1360 498
0 1 16 0 0 12432 0 0 16 30 0 6
1284 225
1284 328
1383 328
1383 508
1366 508
1366 498
1 10 13 0 0 0 0 20 35 0 0 3
1292 661
1292 695
1184 695
11 9 17 0 0 8320 0 34 35 0 0 6
1183 521
1188 521
1188 737
1112 737
1112 722
1120 722
1 10 14 0 0 8320 0 21 34 0 0 3
1292 501
1292 530
1183 530
10 1 15 0 0 4224 0 33 22 0 0 3
1186 379
1288 379
1288 361
10 1 16 0 0 0 0 32 23 0 0 3
1180 225
1284 225
1284 205
11 9 18 0 0 8320 0 33 34 0 0 6
1186 370
1195 370
1195 572
1111 572
1111 557
1119 557
11 9 19 0 0 8320 0 32 33 0 0 6
1180 216
1190 216
1190 421
1114 421
1114 406
1122 406
0 4 4 0 0 0 0 0 18 11 0 5
573 669
575 669
575 558
391 558
391 515
1 3 6 0 0 12288 0 5 18 0 0 5
565 597
575 597
575 552
397 552
397 515
0 2 8 0 0 8192 0 0 18 48 0 4
567 536
567 546
403 546
403 515
0 1 9 0 0 8192 0 0 18 49 0 4
569 480
569 523
409 523
409 515
1 4 20 0 0 4096 0 8 19 0 0 5
565 401
388 401
388 298
387 298
387 231
0 3 21 0 0 8192 0 0 19 42 0 4
582 342
582 287
393 287
393 231
0 2 22 0 0 4096 0 0 19 43 0 3
564 280
399 280
399 231
1 1 23 0 0 12288 0 11 19 0 0 5
563 214
564 214
564 242
405 242
405 231
1 4 20 0 0 8320 0 8 35 0 0 5
565 401
565 465
1015 465
1015 677
1120 677
1 4 21 0 0 4224 0 9 34 0 0 4
563 342
1110 342
1110 512
1119 512
1 4 22 0 0 8320 0 10 33 0 0 5
564 269
564 319
1092 319
1092 361
1122 361
1 4 23 0 0 12416 0 11 32 0 0 6
563 214
564 214
564 181
1075 181
1075 207
1116 207
3 8 24 0 0 4224 0 27 34 0 0 4
1007 547
1110 547
1110 548
1119 548
3 8 25 0 0 4224 0 29 32 0 0 4
995 242
1080 242
1080 243
1116 243
1 1 6 0 0 12416 0 5 15 0 0 6
565 597
589 597
589 560
786 560
786 586
803 586
1 1 8 0 0 12416 0 6 30 0 0 6
564 536
591 536
591 399
783 399
783 432
791 432
1 1 9 0 0 8320 0 7 31 0 0 6
563 480
617 480
617 249
778 249
778 285
785 285
3 8 26 0 0 4224 0 26 35 0 0 4
1012 712
1096 712
1096 713
1120 713
3 8 27 0 0 4224 0 28 33 0 0 2
1002 397
1122 397
2 3 28 0 0 4224 0 26 43 0 0 4
966 721
901 721
901 757
893 757
1 3 29 0 0 4224 0 26 42 0 0 4
966 703
903 703
903 683
895 683
2 3 30 0 0 4224 0 27 41 0 0 4
961 556
904 556
904 595
896 595
1 3 31 0 0 4224 0 27 40 0 0 4
961 538
902 538
902 520
894 520
2 3 32 0 0 4224 0 28 39 0 0 4
956 406
897 406
897 441
889 441
1 3 33 0 0 4224 0 28 38 0 0 4
956 388
895 388
895 367
887 367
3 1 34 0 0 4224 0 36 29 0 0 4
887 210
940 210
940 233
949 233
3 2 35 0 0 4224 0 37 29 0 0 4
885 294
940 294
940 251
949 251
2 0 3 0 0 0 0 41 0 0 0 2
851 604
830 604
1 9 36 0 0 4224 0 3 32 0 0 4
561 157
1070 157
1070 252
1116 252
27
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
384 418 419 441
397 428 405 443
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
379 131 414 154
392 141 400 156
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1296 199 1344 222
1309 209 1330 224
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1098 742 1209 765
1111 752 1195 767
12 Full Adder 4
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1096 570 1207 593
1109 580 1193 595
12 Full Adder 3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1100 421 1209 444
1112 431 1196 446
12 Full Adder 2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1096 264 1205 287
1108 274 1192 289
12 Full Adder 1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1081 710 1120 733
1093 720 1107 735
2 Y3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1077 545 1118 568
1090 555 1104 570
2 Y2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1076 394 1117 417
1089 404 1103 419
2 Y1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1085 216 1124 239
1097 226 1111 241
2 Y0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
473 392 512 415
485 402 499 417
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 322 512 345
484 332 498 347
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 258 510 281
483 268 497 283
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
470 193 509 216
482 203 496 218
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
475 462 516 485
488 472 502 487
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
477 523 518 546
490 533 504 548
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 580 518 603
491 590 505 605
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 657 518 680
491 667 505 682
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
461 141 509 164
474 151 495 166
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1083 649 1124 672
1096 659 1110 674
2 X3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1076 499 1115 522
1088 509 1102 524
2 X2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1077 357 1118 380
1090 367 1104 382
2 X1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
1084 189 1123 212
1096 199 1110 214
2 X0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
944 1452 985 1475
957 1462 971 1477
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
880 1459 919 1482
892 1469 906 1484
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 17
1218 128 1364 151
1231 138 1350 153
17 Arithmetic Output
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
