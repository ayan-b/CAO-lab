CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
170 110 30 90 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
79
13 Logic Switch~
5 765 1574 0 1 11
0 18
0
0 0 21360 90
2 0V
14 0 28 8
3 V14
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3244 0 0
2
43336 0
0
13 Logic Switch~
5 668 1572 0 10 11
0 8 0 0 0 0 0 0 0 0
1
0
0 0 21360 90
2 5V
14 0 28 8
3 V13
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7405 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 713 1574 0 1 11
0 19
0
0 0 21360 90
2 0V
14 0 28 8
3 V12
10 -10 31 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6988 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 549 157 0 10 11
0 68 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -17 6 -9
3 V11
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3858 0 0
2
5.89859e-315 0
0
13 Logic Switch~
5 550 669 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
3 V10
-9 -25 12 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3792 0 0
2
43336 0
0
13 Logic Switch~
5 553 597 0 1 11
0 34
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7557 0 0
2
43336 1
0
13 Logic Switch~
5 552 536 0 1 11
0 45
0
0 0 21360 0
2 0V
-8 -16 6 -8
2 V8
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3913 0 0
2
43336 2
0
13 Logic Switch~
5 551 480 0 10 11
0 49 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V7
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
7686 0 0
2
43336 3
0
13 Logic Switch~
5 553 401 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
357 0 0
2
43336 4
0
13 Logic Switch~
5 551 342 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6967 0 0
2
43336 5
0
13 Logic Switch~
5 552 269 0 1 11
0 53
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3263 0 0
2
43336 6
0
13 Logic Switch~
5 551 214 0 1 11
0 59
0
0 0 21360 0
2 0V
-7 -19 7 -11
2 V3
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
9948 0 0
2
43336 7
0
12 Hex Display~
7 1422 521 0 18 19
10 5 2 4 3 0 0 0 0 0
0 0 1 1 1 1 0 1 13
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7982 0 0
2
43336.1 0
0
14 Logic Display~
6 1309 1438 0 1 2
10 6
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8270 0 0
2
43336.1 0
0
5 4049~
219 1187 1167 0 2 22
0 8 13
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U17F
13 -8 41 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 15 0
1 U
7388 0 0
2
43336.1 1
0
5 4081~
219 1201 1219 0 3 22
0 9 13 7
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U22C
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 18 0
1 U
3351 0 0
2
43336.1 0
0
5 4049~
219 1180 797 0 2 22
0 8 14
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U17E
13 -8 41 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 15 0
1 U
3818 0 0
2
43336.1 1
0
5 4081~
219 1194 849 0 3 22
0 10 14 11
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U22B
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 18 0
1 U
3413 0 0
2
43336.1 0
0
5 4049~
219 1166 464 0 2 22
0 8 15
0
0 0 624 270
4 4049
-7 -24 21 -16
4 U17C
13 -8 41 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 15 0
1 U
8628 0 0
2
43336.1 1
0
5 4081~
219 1180 516 0 3 22
0 12 15 73
0
0 0 624 270
4 4081
-7 -24 21 -16
4 U13D
13 -4 41 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 4 11 0
1 U
7669 0 0
2
43336.1 0
0
14 Logic Display~
6 1308 1130 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4710 0 0
2
43336.1 0
0
14 Logic Display~
6 1303 761 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3594 0 0
2
43336.1 0
0
14 Logic Display~
6 1290 418 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5569 0 0
2
43336.1 0
0
4 4008
219 1201 1312 0 14 29
0 74 75 76 33 77 78 79 16 7
3 6 80 81 82
0
0 0 4848 0
4 4008
-14 -60 14 -52
3 U21
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3128 0 0
2
43336.1 0
0
4 4008
219 1196 945 0 14 29
0 83 84 85 44 86 87 88 17 11
4 9 89 90 91
0
0 0 4848 0
4 4008
-14 -60 14 -52
3 U20
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
5222 0 0
2
43336.1 0
0
5 4071~
219 1099 1425 0 3 22
0 27 28 16
0
0 0 624 0
4 4071
-7 -24 21 -16
4 U19A
-6 -25 22 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 17 0
1 U
6289 0 0
2
43336 10
0
5 4049~
219 937 1468 0 2 22
0 23 26
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 15 0
1 U
3201 0 0
2
43336 9
0
5 4081~
219 1003 1393 0 3 22
0 18 23 27
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13C
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 11 0
1 U
388 0 0
2
43336 8
0
5 4081~
219 1008 1477 0 3 22
0 26 19 28
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13B
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 11 0
1 U
8936 0 0
2
43336 7
0
8 3-In OR~
219 1069 1282 0 4 22
0 20 32 31 33
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U14B
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 1 2 8 9 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 2 12 0
1 U
5590 0 0
2
43336 6
0
5 4082~
219 989 1242 0 5 22
0 23 8 25 24 32
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 16 0
1 U
3980 0 0
2
43336 5
0
5 4082~
219 992 1310 0 5 22
0 30 8 19 29 31
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U18A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 16 0
1 U
3232 0 0
2
43336 4
0
5 4049~
219 920 1298 0 2 22
0 23 30
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U17A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 15 0
1 U
3571 0 0
2
43336 3
0
5 4049~
219 872 1246 0 2 22
0 19 25
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 14 0
1 U
3640 0 0
2
43336 2
0
5 4049~
219 872 1274 0 2 22
0 18 24
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 14 0
1 U
9587 0 0
2
43336 1
0
5 4049~
219 923 1325 0 2 22
0 18 29
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 14 0
1 U
5646 0 0
2
43336 0
0
5 4049~
219 897 975 0 2 22
0 18 40
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 14 0
1 U
7185 0 0
2
43336 10
0
5 4049~
219 846 924 0 2 22
0 18 35
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 14 0
1 U
3167 0 0
2
43336 9
0
5 4049~
219 846 896 0 2 22
0 19 36
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U16A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 14 0
1 U
4184 0 0
2
43336 8
0
5 4049~
219 894 948 0 2 22
0 34 41
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11F
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 10 0
1 U
9609 0 0
2
43336 7
0
5 4082~
219 966 960 0 5 22
0 41 8 19 40 42
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 13 0
1 U
3286 0 0
2
43336 6
0
5 4082~
219 963 892 0 5 22
0 34 8 36 35 43
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U15A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 13 0
1 U
4915 0 0
2
43336 5
0
8 3-In OR~
219 1043 932 0 4 22
0 21 43 42 44
0
0 0 624 0
4 4075
-14 -24 14 -16
4 U14A
-6 -25 22 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 12 0
1 U
8380 0 0
2
43336 4
0
5 4081~
219 982 1127 0 3 22
0 37 19 39
0
0 0 624 0
4 4081
-7 -24 21 -16
4 U13A
-15 -25 13 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 11 0
1 U
869 0 0
2
43336 3
0
5 4081~
219 977 1043 0 3 22
0 18 34 38
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 8 0
1 U
3843 0 0
2
43336 2
0
5 4049~
219 911 1118 0 2 22
0 34 37
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11E
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 10 0
1 U
5584 0 0
2
43336 1
0
5 4071~
219 1073 1075 0 3 22
0 38 39 17
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
5282 0 0
2
43336 0
0
5 4071~
219 1036 723 0 3 22
0 47 48 22
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 5 0
1 U
9831 0 0
2
43336 3
0
5 4049~
219 874 766 0 2 22
0 45 46
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11D
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 10 0
1 U
9598 0 0
2
43336 2
0
5 4081~
219 940 691 0 3 22
0 18 45 47
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 8 0
1 U
3862 0 0
2
43336 1
0
5 4081~
219 945 775 0 3 22
0 46 19 48
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U8C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 8 0
1 U
464 0 0
2
43336 0
0
4 4008
219 1184 599 0 14 29
0 92 93 94 57 95 96 97 22 98
2 10 99 100 101
0
0 0 4848 0
4 4008
-14 -60 14 -52
3 U12
-10 -61 11 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3248 0 0
2
43336 0
0
5 4049~
219 881 652 0 2 22
0 18 52
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11C
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 10 0
1 U
6467 0 0
2
43336 6
0
5 4049~
219 830 601 0 2 22
0 18 50
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11B
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 10 0
1 U
3558 0 0
2
43336 5
0
5 4049~
219 830 573 0 2 22
0 19 51
0
0 0 624 0
4 4049
-7 -24 21 -16
4 U11A
-14 -20 14 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 10 0
1 U
9814 0 0
2
43336 4
0
5 4049~
219 878 625 0 2 22
0 45 54
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U4F
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 6 0
1 U
9595 0 0
2
43336 3
0
5 4082~
219 950 637 0 5 22
0 54 8 19 52 55
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10B
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 9 0
1 U
3455 0 0
2
43336 2
0
5 4082~
219 947 569 0 5 22
0 45 8 51 50 56
0
0 0 624 0
4 4082
-7 -24 21 -16
4 U10A
-15 -28 13 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 9 0
1 U
836 0 0
2
43336 1
0
8 3-In OR~
219 1027 609 0 4 22
0 53 56 55 57
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2C
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 11 12 13 10 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 3 2 0
1 U
3509 0 0
2
43336 0
0
5 4049~
219 871 347 0 2 22
0 18 62
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7F
6 -22 27 -14
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 14 15 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
6760 0 0
2
43336 0
0
5 4049~
219 820 296 0 2 22
0 18 60
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7E
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 11 12 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
4270 0 0
2
43336 0
0
5 4049~
219 820 269 0 2 22
0 19 61
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7D
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 9 10 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
8152 0 0
2
43336 0
0
5 4049~
219 868 320 0 2 22
0 49 64
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 7 6 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
3261 0 0
2
43336 0
0
5 4082~
219 940 332 0 5 22
0 64 8 19 62 65
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3B
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 9 10 11 12 13 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 2 4 0
1 U
727 0 0
2
43336 0
0
5 4082~
219 937 264 0 5 22
0 49 8 61 60 66
0
0 0 624 0
4 4082
-7 -24 21 -16
3 U3A
-12 -28 9 -20
0
15 DVDD=14;DGND=7;
61 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o] %M
0
13 type: digital
5 DIP14
22

0 2 3 4 5 1 2 3 4 5
1 9 10 11 12 13 0 0 0 0
0 1 0
65 0 0 0 2 1 4 0
1 U
5620 0 0
2
43336 0
0
8 3-In OR~
219 1017 304 0 4 22
0 59 66 65 63
0
0 0 624 0
4 4075
-14 -24 14 -16
3 U2A
-3 -25 18 -17
0
15 DVDD=14;DGND=7;
53 %D [%14bi %7bi %1i %2i %3i][%14bo %1o %2o %3o %4o] %M
0
12 type:digital
5 DIP14
22

0 3 4 5 6 3 4 5 6 1
2 8 9 11 12 13 10 0 0 0
0 1 0
65 0 0 0 3 1 2 0
1 U
3286 0 0
2
43336 0
0
5 4049~
219 1156 212 0 2 22
0 8 69
0
0 0 624 270
4 4049
-7 -24 21 -16
3 U7B
16 -8 37 0
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 5 4 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 2 3 0
1 U
8481 0 0
2
43336 0
0
5 4081~
219 1170 264 0 3 22
0 68 69 67
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U5C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
8955 0 0
2
43336 0
0
5 4081~
219 924 471 0 3 22
0 70 19 72
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
534 0 0
2
43336 3
0
5 4081~
219 919 387 0 3 22
0 18 49 71
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U5A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
4680 0 0
2
43336 2
0
5 4049~
219 853 462 0 2 22
0 49 70
0
0 0 624 0
4 4049
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
14 DVDD=1;DGND=8;
35 %D [%1bi %8bi %1i][%1bo %1o %2o] %M
0
12 type:digital
5 DIP16
22

0 3 2 3 2 5 4 7 6 9
10 11 12 14 15 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
3540 0 0
2
43336 1
0
5 4071~
219 1015 419 0 3 22
0 71 72 58
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
3974 0 0
2
43336 0
0
14 Logic Display~
6 753 107 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9365 0 0
2
43336 0
0
12 Hex Display~
7 400 491 0 18 19
10 49 45 34 23 0 0 0 0 0
0 1 1 1 1 0 1 1 9
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
369 0 0
2
5.89859e-315 5.3568e-315
0
12 Hex Display~
7 396 207 0 18 19
10 59 53 21 20 0 0 0 0 0
0 1 0 0 1 1 1 0 12
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3927 0 0
2
5.89859e-315 5.36716e-315
0
14 Logic Display~
6 1284 187 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9659 0 0
2
5.89859e-315 5.39824e-315
0
14 Logic Display~
6 719 114 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7205 0 0
2
5.89859e-315 5.40342e-315
0
14 Logic Display~
6 677 118 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3413 0 0
2
5.89859e-315 5.4086e-315
0
4 4008
219 1178 369 0 14 29
0 102 103 104 63 105 106 107 58 67
5 12 108 109 110
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
4708 0 0
2
43336 10
0
138
2 0 2 0 0 8192 0 13 0 0 20 5
1425 545
1425 554
1295 554
1295 541
1290 541
0 4 3 0 0 8320 0 0 13 18 0 3
1308 1170
1413 1170
1413 545
0 3 4 0 0 8320 0 0 13 19 0 3
1303 804
1419 804
1419 545
1 0 5 0 0 12288 0 13 0 0 130 4
1431 545
1431 549
1277 549
1277 378
11 1 6 0 0 8320 0 24 14 0 0 5
1233 1312
1296 1312
1296 1464
1309 1464
1309 1456
3 9 7 0 0 12416 0 16 24 0 0 5
1199 1242
1199 1257
1156 1257
1156 1348
1169 1348
1 0 8 0 0 8192 0 15 0 0 129 3
1190 1149
1190 1145
669 1145
11 1 9 0 0 8320 0 25 16 0 0 5
1228 945
1232 945
1232 1189
1208 1189
1208 1197
1 11 10 0 0 4224 0 18 52 0 0 5
1201 827
1201 649
1224 649
1224 599
1216 599
3 9 11 0 0 12416 0 18 25 0 0 5
1192 872
1192 890
1151 890
1151 981
1164 981
0 0 8 0 0 0 0 0 0 12 129 3
684 825
684 824
669 824
1 0 8 0 0 0 0 17 0 0 0 5
1183 779
1183 780
1152 780
1152 825
681 825
1 0 8 0 0 0 0 19 0 0 129 4
1169 446
1139 446
1139 491
668 491
11 1 12 0 0 8320 0 79 20 0 0 5
1210 369
1214 369
1214 486
1187 486
1187 494
2 2 13 0 0 4224 0 16 15 0 0 2
1190 1197
1190 1185
2 2 14 0 0 4224 0 18 17 0 0 2
1183 827
1183 815
2 2 15 0 0 4224 0 20 19 0 0 2
1169 494
1169 482
10 1 3 0 0 0 0 24 21 0 0 3
1233 1321
1308 1321
1308 1148
10 1 4 0 0 0 0 25 22 0 0 4
1228 954
1228 952
1303 952
1303 779
10 1 2 0 0 12416 0 52 23 0 0 4
1216 608
1216 609
1290 609
1290 436
3 8 16 0 0 8320 0 26 24 0 0 4
1132 1425
1161 1425
1161 1339
1169 1339
3 8 17 0 0 8320 0 47 25 0 0 4
1106 1075
1156 1075
1156 972
1164 972
1 0 18 0 0 4096 0 35 0 0 128 2
857 1274
753 1274
1 0 18 0 0 4096 0 36 0 0 128 4
908 1325
758 1325
758 1326
753 1326
3 0 19 0 0 8192 0 32 0 0 108 3
968 1315
968 1317
717 1317
2 0 8 0 0 0 0 32 0 0 129 3
968 1306
968 1307
669 1307
1 0 19 0 0 0 0 34 0 0 108 2
857 1246
717 1246
2 0 8 0 0 0 0 31 0 0 129 4
965 1238
897 1238
897 1239
669 1239
0 0 19 0 0 0 0 0 0 45 108 2
823 1486
717 1486
0 0 18 0 0 0 0 0 0 46 128 2
870 1384
753 1384
1 0 20 0 0 8320 0 9 0 0 52 5
565 401
622 401
622 1191
810 1191
811 1192
0 0 21 0 0 8192 0 0 0 33 136 3
594 381
582 381
582 342
1 0 21 0 0 12416 0 43 0 0 0 4
1030 923
1030 859
594 859
594 378
1 0 18 0 0 0 0 37 0 0 128 2
882 975
753 975
3 0 19 0 0 0 0 41 0 0 108 3
942 965
942 970
717 970
2 0 8 0 0 0 0 41 0 0 129 3
942 956
942 961
669 961
1 0 18 0 0 0 0 38 0 0 128 2
831 924
753 924
1 0 19 0 0 0 0 39 0 0 108 2
831 896
717 896
2 0 8 0 0 0 0 42 0 0 129 2
939 888
669 888
0 0 18 0 0 0 0 0 0 63 128 2
844 1034
753 1034
3 8 22 0 0 8320 0 48 52 0 0 4
1069 723
1144 723
1144 626
1152 626
0 0 23 0 0 4096 0 0 0 53 47 3
842 1229
842 1430
914 1430
2 4 24 0 0 8320 0 35 31 0 0 3
893 1274
893 1256
965 1256
2 3 25 0 0 4224 0 34 31 0 0 4
893 1246
957 1246
957 1247
965 1247
2 0 19 0 0 0 0 29 0 0 0 2
984 1486
820 1486
1 0 18 0 0 0 0 28 0 0 30 2
979 1384
867 1384
1 2 23 0 0 0 0 27 28 0 0 4
922 1468
914 1468
914 1402
979 1402
1 2 26 0 0 4224 0 29 27 0 0 2
984 1468
958 1468
3 1 27 0 0 4224 0 28 26 0 0 4
1024 1393
1077 1393
1077 1416
1086 1416
3 2 28 0 0 4224 0 29 26 0 0 4
1029 1477
1077 1477
1077 1434
1086 1434
4 2 29 0 0 4224 0 32 36 0 0 4
968 1324
952 1324
952 1325
944 1325
0 1 20 0 0 0 0 0 30 31 0 4
811 1192
1048 1192
1048 1273
1056 1273
0 1 23 0 0 12416 0 0 31 131 0 5
579 669
579 674
585 674
585 1229
965 1229
1 0 23 0 0 0 0 33 0 0 53 3
905 1298
901 1298
901 1229
2 1 30 0 0 4224 0 33 32 0 0 4
941 1298
960 1298
960 1297
968 1297
3 5 31 0 0 4224 0 30 32 0 0 4
1056 1291
1021 1291
1021 1310
1013 1310
2 5 32 0 0 8320 0 30 31 0 0 4
1057 1282
1018 1282
1018 1242
1010 1242
4 4 33 0 0 12416 0 30 24 0 0 4
1102 1282
1120 1282
1120 1303
1169 1303
0 0 34 0 0 4096 0 0 0 69 64 3
816 879
816 1080
888 1080
2 4 35 0 0 8320 0 38 42 0 0 3
867 924
867 906
939 906
2 3 36 0 0 4224 0 39 42 0 0 4
867 896
931 896
931 897
939 897
2 0 19 0 0 0 0 44 0 0 108 2
958 1136
717 1136
1 0 18 0 0 0 0 45 0 0 40 2
953 1034
841 1034
1 2 34 0 0 0 0 46 45 0 0 4
896 1118
888 1118
888 1052
953 1052
1 2 37 0 0 4224 0 44 46 0 0 2
958 1118
932 1118
3 1 38 0 0 4224 0 45 47 0 0 4
998 1043
1051 1043
1051 1066
1060 1066
3 2 39 0 0 4224 0 44 47 0 0 4
1003 1127
1051 1127
1051 1084
1060 1084
4 2 40 0 0 4224 0 41 37 0 0 4
942 974
926 974
926 975
918 975
0 1 34 0 0 8320 0 0 42 132 0 3
574 597
574 879
939 879
1 0 34 0 0 0 0 40 0 0 69 3
879 948
875 948
875 879
2 1 41 0 0 4224 0 40 41 0 0 4
915 948
934 948
934 947
942 947
3 5 42 0 0 4224 0 43 41 0 0 4
1030 941
995 941
995 960
987 960
2 5 43 0 0 8320 0 43 42 0 0 4
1031 932
992 932
992 892
984 892
4 4 44 0 0 12416 0 43 25 0 0 4
1076 932
1094 932
1094 936
1164 936
1 0 45 0 0 8192 0 56 0 0 78 4
863 625
829 625
829 732
851 732
2 0 19 0 0 0 0 51 0 0 108 2
921 784
718 784
1 0 18 0 0 0 0 50 0 0 128 4
916 682
804 682
804 683
753 683
1 2 45 0 0 0 0 49 50 0 0 4
859 766
851 766
851 700
916 700
1 2 46 0 0 4224 0 51 49 0 0 2
921 766
895 766
3 1 47 0 0 4224 0 50 48 0 0 4
961 691
1014 691
1014 714
1023 714
3 2 48 0 0 4224 0 51 48 0 0 4
966 775
1014 775
1014 732
1023 732
1 0 18 0 0 0 0 53 0 0 128 2
866 652
753 652
3 0 19 0 0 0 0 57 0 0 108 3
926 642
926 640
717 640
2 0 8 0 0 0 0 57 0 0 129 3
926 633
926 632
668 632
1 0 18 0 0 0 0 54 0 0 128 2
815 601
753 601
1 0 19 0 0 0 0 55 0 0 108 2
815 573
717 573
2 0 8 0 0 0 0 58 0 0 129 2
923 565
668 565
0 0 49 0 0 8192 0 0 0 124 116 3
830 434
772 434
772 251
2 4 50 0 0 8320 0 54 58 0 0 3
851 601
851 583
923 583
2 3 51 0 0 4224 0 55 58 0 0 4
851 573
915 573
915 574
923 574
4 2 52 0 0 4224 0 57 53 0 0 4
926 651
910 651
910 652
902 652
1 1 53 0 0 12416 0 11 59 0 0 6
564 269
640 269
640 519
1006 519
1006 600
1014 600
1 1 45 0 0 16512 0 7 58 0 0 5
564 536
564 538
586 538
586 556
923 556
1 0 45 0 0 0 0 56 0 0 93 3
863 625
859 625
859 556
2 1 54 0 0 4224 0 56 57 0 0 4
899 625
918 625
918 624
926 624
3 5 55 0 0 4224 0 59 57 0 0 4
1014 618
979 618
979 637
971 637
2 5 56 0 0 8320 0 59 58 0 0 4
1015 609
976 609
976 569
968 569
4 4 57 0 0 12416 0 59 52 0 0 4
1060 609
1078 609
1078 590
1152 590
1 0 18 0 0 0 0 70 0 0 128 2
895 378
753 378
3 8 58 0 0 4224 0 72 79 0 0 4
1048 419
1138 419
1138 396
1146 396
2 0 8 0 0 0 0 64 0 0 129 3
916 328
916 334
668 334
3 0 19 0 0 0 0 64 0 0 108 3
916 337
916 339
717 339
1 0 18 0 0 0 0 60 0 0 128 2
856 347
753 347
1 0 18 0 0 0 0 61 0 0 128 2
805 296
753 296
1 0 19 0 0 0 0 62 0 0 108 2
805 269
717 269
2 0 8 0 0 0 0 65 0 0 129 4
913 260
845 260
845 259
668 259
1 1 59 0 0 16512 0 66 12 0 0 5
1004 295
1004 215
855 215
855 214
563 214
1 1 19 0 0 16528 0 3 77 0 0 11
714 1561
716 1561
716 1491
717 1491
717 789
718 789
718 645
717 645
717 139
719 139
719 132
0 1 8 0 0 0 0 0 67 129 0 3
672 187
1159 187
1159 194
2 4 60 0 0 4224 0 61 65 0 0 4
841 296
905 296
905 278
913 278
3 2 61 0 0 4224 0 65 62 0 0 2
913 269
841 269
4 2 62 0 0 4224 0 64 60 0 0 4
916 346
900 346
900 347
892 347
0 4 63 0 0 4224 0 0 79 120 0 4
1062 304
1138 304
1138 360
1146 360
1 0 49 0 0 0 0 63 0 0 116 3
853 320
849 320
849 251
2 1 64 0 0 4224 0 63 64 0 0 4
889 320
908 320
908 319
916 319
0 1 49 0 0 12416 0 0 65 134 0 4
567 480
603 480
603 251
913 251
3 5 65 0 0 4224 0 66 64 0 0 4
1004 313
969 313
969 332
961 332
2 5 66 0 0 8320 0 66 65 0 0 4
1005 304
966 304
966 264
958 264
9 3 67 0 0 8320 0 79 68 0 0 5
1146 405
1142 405
1142 295
1168 295
1168 287
4 0 63 0 0 0 0 66 0 0 0 2
1050 304
1068 304
1 1 68 0 0 4224 0 4 68 0 0 3
561 157
1177 157
1177 242
2 2 69 0 0 4224 0 68 67 0 0 2
1159 242
1159 230
2 0 19 0 0 0 0 69 0 0 108 2
900 480
717 480
1 2 49 0 0 0 0 71 70 0 0 4
838 462
830 462
830 396
895 396
1 2 70 0 0 4224 0 69 71 0 0 2
900 462
874 462
3 1 71 0 0 4224 0 70 72 0 0 4
940 387
993 387
993 410
1002 410
3 2 72 0 0 4224 0 69 72 0 0 4
945 471
993 471
993 428
1002 428
1 1 18 0 0 16512 0 73 1 0 0 6
753 125
752 125
752 266
753 266
753 1561
766 1561
1 1 8 0 0 24704 0 78 2 0 0 7
677 136
672 136
672 192
668 192
668 632
669 632
669 1559
10 1 5 0 0 8320 0 79 76 0 0 3
1210 378
1284 378
1284 205
1 4 23 0 0 0 0 5 74 0 0 5
562 669
580 669
580 558
391 558
391 515
1 3 34 0 0 0 0 6 74 0 0 5
565 597
575 597
575 552
397 552
397 515
0 2 45 0 0 0 0 0 74 93 0 4
567 538
567 546
403 546
403 515
1 1 49 0 0 0 0 8 74 0 0 5
563 480
569 480
569 523
409 523
409 515
1 4 20 0 0 0 0 9 75 0 0 5
565 401
388 401
388 298
387 298
387 231
1 3 21 0 0 0 0 10 75 0 0 5
563 342
582 342
582 287
393 287
393 231
1 2 53 0 0 0 0 11 75 0 0 7
564 269
573 269
573 279
564 279
564 280
399 280
399 231
1 1 59 0 0 0 0 12 75 0 0 5
563 214
564 214
564 242
405 242
405 231
17
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 34
856 1596 1083 1620
867 1605 1071 1621
34 ARITHMETIC LOGIC UNIT (METHOD III)
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 12
1227 129 1340 144
1241 140 1325 151
12 Final Output
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
654 1588 693 1611
666 1598 680 1613
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
704 1590 745 1613
717 1600 731 1615
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
763 1590 802 1613
775 1600 789 1615
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
461 141 509 164
474 151 495 166
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 657 518 680
491 667 505 682
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
479 580 518 603
491 590 505 605
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
477 523 518 546
490 533 504 548
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
475 462 516 485
488 472 502 487
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
470 193 509 216
482 203 496 218
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 258 510 281
483 268 497 283
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
471 322 512 345
484 332 498 347
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
473 392 512 415
485 402 499 417
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
1296 199 1344 222
1309 209 1330 224
3 LSB
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
379 131 414 154
392 141 400 156
1 A
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
384 418 419 441
397 428 405 443
1 B
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
