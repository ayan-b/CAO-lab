CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
30 380 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
41
13 Logic Switch~
5 314 145 0 1 11
0 13
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3165 0 0
2
43340.6 0
0
13 Logic Switch~
5 317 218 0 1 11
0 12
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7874 0 0
2
43340.6 1
0
13 Logic Switch~
5 323 294 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3280 0 0
2
43340.6 2
0
13 Logic Switch~
5 326 380 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3122 0 0
2
43340.6 3
0
13 Logic Switch~
5 330 470 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
6242 0 0
2
43340.6 4
0
13 Logic Switch~
5 333 544 0 1 11
0 8
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8862 0 0
2
43340.6 5
0
13 Logic Switch~
5 316 71 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V7
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3202 0 0
2
43340.6 6
0
13 Logic Switch~
5 374 637 0 1 11
0 14
0
0 0 21360 90
2 0V
11 0 25 8
2 V8
11 -10 25 -2
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5657 0 0
2
43340.6 7
0
7 Ground~
168 889 198 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3554 0 0
2
5.8986e-315 0
0
12 Hex Display~
7 898 170 0 16 19
10 7 6 5 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4316 0 0
2
43340.6 8
0
7 Ground~
168 205 496 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3739 0 0
2
43340.6 9
0
12 Hex Display~
7 229 450 0 16 19
10 10 9 8 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
7606 0 0
2
43340.6 10
0
7 Ground~
168 187 195 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3741 0 0
2
43340.6 11
0
12 Hex Display~
7 221 159 0 16 19
10 13 12 11 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
369 0 0
2
43340.6 12
0
5 4071~
219 645 539 0 3 22
0 20 23 17
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U9A
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
8773 0 0
2
43340.6 13
0
5 4069~
219 522 607 0 2 22
0 3 4
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 2 5 0
1 U
7981 0 0
2
43340.6 14
0
5 4069~
219 513 510 0 2 22
0 8 21
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U8A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 5 0
1 U
4205 0 0
2
43340.6 15
0
5 4081~
219 602 598 0 3 22
0 8 4 23
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2D
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
3375 0 0
2
43340.6 16
0
5 4081~
219 597 501 0 3 22
0 21 14 20
0
0 0 624 692
4 4081
-7 -24 21 -16
3 U2C
-14 -25 7 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
719 0 0
2
43340.6 17
0
5 4071~
219 638 326 0 3 22
0 18 25 22
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1D
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3749 0 0
2
43340.6 18
0
5 4069~
219 501 389 0 2 22
0 3 24
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7F
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 13 12 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 6 3 0
1 U
3871 0 0
2
43340.6 19
0
5 4069~
219 494 295 0 2 22
0 9 19
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7E
-11 -22 10 -14
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 11 10 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 5 3 0
1 U
4393 0 0
2
43340.6 20
0
5 4081~
219 590 380 0 3 22
0 9 24 25
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U2B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
6229 0 0
2
43340.6 21
0
5 4081~
219 581 286 0 3 22
0 19 14 18
0
0 0 624 692
4 4081
-7 -24 21 -16
3 U2A
-14 -25 7 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3757 0 0
2
43340.6 22
0
5 4081~
219 601 2752 0 3 22
0 30 37 29
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6A
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 1 2 0
1 U
352 0 0
2
43340.6 23
0
5 4081~
219 602 2849 0 3 22
0 26 27 28
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6B
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
3372 0 0
2
43340.6 24
0
5 4069~
219 511 2743 0 2 22
0 26 30
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7A
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 1 2 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 1 3 0
1 U
4911 0 0
2
43340.6 25
0
5 4069~
219 519 2858 0 2 22
0 38 27
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7B
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 3 4 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 512 6 2 3 0
1 U
7574 0 0
2
43340.6 26
0
5 4071~
219 676 2793 0 3 22
0 29 28 39
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1B
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 512 4 2 1 0
1 U
6601 0 0
2
43340.6 27
0
14 Logic Display~
6 827 564 0 1 2
10 32
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8531 0 0
2
43340.6 28
0
14 Logic Display~
6 825 477 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6532 0 0
2
43340.6 29
0
14 Logic Display~
6 814 297 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3621 0 0
2
43340.6 30
0
14 Logic Display~
6 808 91 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5174 0 0
2
43340.6 31
0
4 4008
219 729 156 0 14 29
0 40 41 42 13 43 44 45 31 3
7 34 46 47 48
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U3
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
5452 0 0
2
43340.6 32
0
4 4008
219 735 333 0 14 29
0 49 50 51 12 52 53 54 22 34
6 33 55 56 57
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U4
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3626 0 0
2
43340.6 33
0
4 4008
219 736 519 0 14 29
0 58 59 60 11 61 62 63 17 33
5 32 64 65 66
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U5
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3806 0 0
2
43340.6 34
0
5 4071~
219 637 129 0 3 22
0 16 36 31
0
0 0 624 0
4 4071
-7 -24 21 -16
3 U1C
-3 -25 18 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3389 0 0
2
43340.6 35
0
5 4069~
219 488 175 0 2 22
0 3 35
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7C
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 5 6 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 3 3 0
1 U
9156 0 0
2
43340.6 36
0
5 4069~
219 481 95 0 2 22
0 10 15
0
0 0 624 0
4 4069
-7 -24 21 -16
3 U7D
-11 -20 10 -12
0
15 DVDD=14;DGND=7;
37 %D [%14bi %7bi %1i][%14bo %1o %2o] %M
0
12 type:digital
5 DIP14
22

0 9 8 1 2 3 4 5 6 9
8 11 10 13 12 0 0 0 0 0
0 1 0
65 0 0 0 6 4 3 0
1 U
5810 0 0
2
43340.6 37
0
5 4081~
219 568 167 0 3 22
0 10 35 36
0
0 0 624 0
4 4081
-7 -24 21 -16
3 U6C
-12 -25 9 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
8260 0 0
2
43340.6 38
0
5 4081~
219 564 87 0 3 22
0 15 14 16
0
0 0 624 692
4 4081
-7 -24 21 -16
3 U6D
-14 -25 7 -17
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
7286 0 0
2
43340.6 39
0
54
1 4 2 0 0 4096 0 9 10 0 0 2
889 192
889 194
1 0 3 0 0 8192 0 16 0 0 3 3
507 607
421 607
421 388
0 1 3 0 0 0 0 0 21 47 0 3
421 192
421 389
486 389
2 2 4 0 0 4224 0 18 16 0 0 2
578 607
543 607
0 3 5 0 0 8320 0 0 10 44 0 3
825 528
895 528
895 194
2 0 6 0 0 4224 0 10 0 0 45 3
901 194
901 342
814 342
0 1 7 0 0 8320 0 0 10 46 0 4
808 165
808 202
907 202
907 194
1 4 2 0 0 8192 0 11 12 0 0 4
205 490
205 482
220 482
220 474
1 3 8 0 0 12288 0 6 12 0 0 5
345 544
360 544
360 492
226 492
226 474
1 2 9 0 0 12288 0 5 12 0 0 5
342 470
351 470
351 487
232 487
232 474
1 1 10 0 0 12288 0 4 12 0 0 5
338 380
403 380
403 482
238 482
238 474
4 1 2 0 0 8320 0 14 13 0 0 4
212 183
212 181
187 181
187 189
1 3 11 0 0 12288 0 3 14 0 0 5
335 294
340 294
340 201
218 201
218 183
1 2 12 0 0 12288 0 2 14 0 0 5
329 218
334 218
334 196
224 196
224 183
1 1 13 0 0 12288 0 1 14 0 0 5
326 145
331 145
331 191
230 191
230 183
1 2 14 0 0 12416 0 8 41 0 0 5
375 624
375 492
376 492
376 78
540 78
2 1 15 0 0 8320 0 39 41 0 0 3
502 95
502 96
540 96
3 1 16 0 0 8320 0 41 37 0 0 4
585 87
614 87
614 120
624 120
8 3 17 0 0 12416 0 36 15 0 0 4
704 546
700 546
700 539
678 539
0 2 14 0 0 0 0 0 24 16 0 2
376 277
557 277
3 1 18 0 0 8320 0 24 20 0 0 4
602 286
614 286
614 317
625 317
2 1 19 0 0 4224 0 22 24 0 0 2
515 295
557 295
2 0 14 0 0 0 0 19 0 0 16 2
573 492
376 492
3 1 20 0 0 8320 0 19 15 0 0 4
618 501
623 501
623 530
632 530
2 1 21 0 0 4224 0 17 19 0 0 2
534 510
573 510
0 1 8 0 0 0 0 0 6 30 0 2
434 544
345 544
0 1 9 0 0 8320 0 0 5 32 0 4
428 328
351 328
351 470
342 470
8 3 22 0 0 8320 0 35 20 0 0 4
703 360
683 360
683 326
671 326
1 4 11 0 0 12416 0 3 36 0 0 6
335 294
358 294
358 414
661 414
661 510
704 510
1 1 8 0 0 12416 0 17 18 0 0 4
498 510
434 510
434 589
578 589
3 2 23 0 0 8320 0 18 15 0 0 4
623 598
625 598
625 548
632 548
1 1 9 0 0 0 0 22 23 0 0 4
479 295
428 295
428 371
566 371
2 2 24 0 0 4224 0 23 21 0 0 2
566 389
522 389
3 2 25 0 0 8320 0 23 20 0 0 4
611 380
616 380
616 335
625 335
1 1 26 0 0 8320 0 27 26 0 0 4
496 2743
492 2743
492 2840
578 2840
2 2 27 0 0 4224 0 26 28 0 0 2
578 2858
540 2858
3 2 28 0 0 8320 0 26 29 0 0 4
623 2849
632 2849
632 2802
663 2802
1 3 29 0 0 4224 0 29 25 0 0 4
663 2784
630 2784
630 2752
622 2752
1 2 30 0 0 4224 0 25 27 0 0 2
577 2743
532 2743
8 3 31 0 0 8320 0 34 37 0 0 4
697 183
686 183
686 129
670 129
11 1 32 0 0 8320 0 36 30 0 0 5
768 519
779 519
779 608
827 608
827 582
11 9 33 0 0 8320 0 35 36 0 0 6
767 333
791 333
791 579
682 579
682 555
704 555
11 9 34 0 0 8320 0 34 35 0 0 5
761 156
778 156
778 391
703 391
703 369
10 1 5 0 0 0 0 36 31 0 0 3
768 528
825 528
825 495
10 1 6 0 0 0 0 35 32 0 0 3
767 342
814 342
814 315
10 1 7 0 0 0 0 34 33 0 0 3
761 165
808 165
808 109
0 9 3 0 0 8320 0 0 34 48 0 3
421 175
421 192
697 192
1 1 3 0 0 0 0 38 7 0 0 4
473 175
337 175
337 71
328 71
1 0 10 0 0 8320 0 4 0 0 51 4
338 380
403 380
403 117
421 117
2 2 35 0 0 4224 0 40 38 0 0 4
544 176
507 176
507 175
509 175
1 1 10 0 0 0 0 39 40 0 0 4
466 95
421 95
421 158
544 158
3 2 36 0 0 8320 0 40 37 0 0 4
589 167
615 167
615 138
624 138
1 4 12 0 0 4224 0 2 35 0 0 4
329 218
696 218
696 324
703 324
1 4 13 0 0 8336 0 1 34 0 0 4
326 145
326 146
697 146
697 147
9
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
361 646 390 670
372 654 378 670
1 S
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 3
256 65 301 89
266 73 290 89
3 Cin
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
264 130 301 154
274 138 290 154
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
267 204 304 228
277 212 293 228
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
269 282 306 306
279 290 295 306
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
270 368 307 392
280 376 296 392
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
273 457 310 481
283 465 299 481
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
273 531 310 555
283 539 299 555
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 49
415 676 732 700
426 684 720 700
49 ARITHMETIC LOGIC UNIT (acc. to given truth table)
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
