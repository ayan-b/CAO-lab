CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 80 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
10 G:\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
36
13 Logic Switch~
5 124 129 0 1 11
0 24
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V9
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89858e-315 0
0
13 Logic Switch~
5 794 440 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-8 -16 6 -8
3 V15
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
391 0 0
2
5.89858e-315 5.26354e-315
0
13 Logic Switch~
5 1120 594 0 1 11
0 14
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V14
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
5.89858e-315 5.30499e-315
0
13 Logic Switch~
5 1146 14 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V13
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
5.89858e-315 5.32571e-315
0
13 Logic Switch~
5 622 27 0 1 11
0 9
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V12
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
5.89858e-315 5.34643e-315
0
13 Logic Switch~
5 304 16 0 1 11
0 25
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V8
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
5.89858e-315 5.3568e-315
0
13 Logic Switch~
5 341 370 0 1 11
0 26
0
0 0 21360 0
2 0V
-6 -16 8 -8
3 V11
-10 -26 11 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8901 0 0
2
5.89858e-315 5.36716e-315
0
13 Logic Switch~
5 304 115 0 10 11
0 23 0 0 0 0 0 0 0 0
1
0
0 0 20848 0
2 5V
-2 -12 12 -4
2 V1
-2 -22 12 -14
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
7361 0 0
2
5.89858e-315 5.37752e-315
0
13 Logic Switch~
5 302 92 0 1 11
0 22
0
0 0 21360 0
2 0V
-7 -15 7 -7
2 V7
-6 -25 8 -17
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
4747 0 0
2
5.89858e-315 5.38788e-315
0
13 Logic Switch~
5 306 52 0 10 11
0 21 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
972 0 0
2
5.89858e-315 5.39306e-315
0
13 Logic Switch~
5 52 122 0 10 11
0 20 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V5
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3472 0 0
2
5.89858e-315 5.39824e-315
0
13 Logic Switch~
5 116 321 0 1 11
0 30
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
9998 0 0
2
5.89858e-315 5.40342e-315
0
13 Logic Switch~
5 118 258 0 10 11
0 31 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3536 0 0
2
5.89858e-315 5.4086e-315
0
13 Logic Switch~
5 118 194 0 10 11
0 32 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -27 8 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
4597 0 0
2
5.89858e-315 5.41378e-315
0
9 2-In XOR~
219 1110 260 0 3 22
0 7 5 17
0
0 0 624 0
5 74F86
-18 -24 17 -16
3 U6A
-5 -25 16 -17
0
15 DVCC=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 4 5 6
9 10 8 12 13 11 0 0 0 0
0 6 0
65 0 0 0 4 1 4 0
1 U
3835 0 0
2
5.89858e-315 5.41896e-315
0
14 Logic Display~
6 1300 172 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
5.89858e-315 5.42414e-315
0
5 4013~
219 1211 206 0 6 22
0 4 8 13 4 33 15
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 5 0
1 U
5616 0 0
2
5.89858e-315 5.42933e-315
0
14 Logic Display~
6 1303 318 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9323 0 0
2
5.89858e-315 5.43192e-315
0
14 Logic Display~
6 1297 25 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
5.89858e-315 5.43451e-315
0
5 4013~
219 1176 85 0 6 22
0 4 7 13 4 34 16
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U7A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 5 0
1 U
3108 0 0
2
5.89858e-315 5.4371e-315
0
5 4013~
219 1246 373 0 6 22
0 4 17 13 4 35 10
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5B
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 8 9 11 10 12 13 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 2 3 0
1 U
4299 0 0
2
5.89858e-315 5.43969e-315
0
5 4013~
219 1074 486 0 6 22
0 4 18 13 14 36 11
0
0 0 4720 0
4 4013
10 -60 38 -52
3 U5A
22 -61 43 -53
0
15 DVDD=14;DGND=7;
65 %D [%14bi %7bi %1i %2i %3i %4i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 6 5 3 4 2 1 6 5 3
4 2 1 8 9 11 10 12 13 0
0 9 0
65 0 0 512 2 1 3 0
1 U
9672 0 0
2
5.89858e-315 5.44228e-315
0
14 Logic Display~
6 1304 417 0 1 2
10 11
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7876 0 0
2
5.89858e-315 5.44487e-315
0
5 7425~
219 936 458 0 6 22
0 8 3 19 2 12 18
0
0 0 624 0
4 7425
-14 -24 14 -16
3 U4A
-3 19 18 27
0
15 DVCC=14;DGND=7;
69 %D [%14bi %7bi %1i %2i %3i %4i %5i][%14bo %1o %2o %3o %4o %5o %6o] %M
0
12 type:digital
5 DIP14
22

0 5 4 2 1 3 6 5 4 2
1 3 6 9 10 12 13 11 8 0
0 6 0
65 0 0 0 2 1 2 0
1 U
6369 0 0
2
5.89858e-315 5.44746e-315
0
14 Logic Display~
6 968 37 0 1 2
10 7
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9172 0 0
2
5.89858e-315 5.45005e-315
0
14 Logic Display~
6 980 323 0 1 2
10 3
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7100 0 0
2
5.89858e-315 5.45264e-315
0
14 Logic Display~
6 978 263 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3820 0 0
2
5.89858e-315 5.45523e-315
0
14 Logic Display~
6 972 210 0 1 2
10 19
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7678 0 0
2
5.89858e-315 5.45782e-315
0
14 Logic Display~
6 971 151 0 1 2
10 8
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
961 0 0
2
5.89858e-315 5.46041e-315
0
5 4030~
219 589 215 0 3 22
0 24 20 6
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3D
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 1 0
1 U
3178 0 0
2
5.89858e-315 0
0
5 4030~
219 226 310 0 3 22
0 30 20 28
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3C
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 1 0
1 U
3409 0 0
2
5.89858e-315 5.26354e-315
0
5 4030~
219 226 259 0 3 22
0 31 20 29
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3B
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 1 0
1 U
3951 0 0
2
5.89858e-315 5.30499e-315
0
5 4030~
219 226 207 0 3 22
0 32 20 27
0
0 0 624 0
4 4030
-7 -24 21 -16
3 U3A
-5 -25 16 -17
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 1 0
1 U
8885 0 0
2
5.89858e-315 5.32571e-315
0
7 Pulser~
4 132 539 0 10 12
0 37 38 13 39 0 0 5 5 1
7
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
3780 0 0
2
5.89858e-315 5.34643e-315
0
4 4008
219 820 189 0 14 29
0 9 9 9 25 9 9 9 6 5
8 7 40 41 42
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U2
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9265 0 0
2
5.89858e-315 5.3568e-315
0
4 4008
219 485 250 0 14 29
0 26 21 22 23 26 27 29 28 20
3 2 19 5 43
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
9442 0 0
2
5.89858e-315 5.36716e-315
0
58
0 4 2 0 0 4096 0 0 24 4 0 3
884 290
884 472
919 472
2 0 3 0 0 8192 0 24 0 0 3 5
919 454
915 454
915 354
964 354
964 349
10 1 3 0 0 4224 0 36 26 0 0 5
517 259
961 259
961 349
980 349
980 341
1 11 2 0 0 8320 0 27 36 0 0 5
978 281
978 290
671 290
671 250
517 250
4 0 4 0 0 8192 0 21 0 0 25 3
1246 379
1246 409
1074 409
0 2 5 0 0 8320 0 0 15 7 0 5
742 225
742 394
1086 394
1086 269
1094 269
9 13 5 0 0 0 0 35 36 0 0 6
788 225
626 225
626 233
525 233
525 232
517 232
8 3 6 0 0 12416 0 35 30 0 0 4
788 216
773 216
773 215
622 215
1 0 7 0 0 8320 0 15 0 0 10 3
1094 251
1064 251
1064 59
1 2 7 0 0 0 0 25 20 0 0 5
968 55
968 59
1144 59
1144 49
1152 49
1 2 8 0 0 8320 0 29 17 0 0 5
971 169
971 173
1179 173
1179 170
1187 170
7 0 9 0 0 8192 0 35 0 0 13 3
788 207
788 198
778 198
6 0 9 0 0 4096 0 35 0 0 14 3
788 198
777 198
777 189
5 0 9 0 0 8320 0 35 0 0 17 3
788 189
690 189
690 27
0 3 9 0 0 0 0 0 35 16 0 3
783 162
783 171
788 171
0 2 9 0 0 0 0 0 35 17 0 3
780 152
780 162
788 162
1 1 9 0 0 0 0 5 35 0 0 4
634 27
780 27
780 153
788 153
6 1 10 0 0 12416 0 21 18 0 0 5
1270 337
1286 337
1286 344
1303 344
1303 336
1 6 11 0 0 8320 0 23 22 0 0 5
1304 435
1304 462
1112 462
1112 450
1098 450
1 5 12 0 0 8320 0 2 24 0 0 6
806 440
806 430
941 430
941 429
941 429
941 437
3 0 13 0 0 4096 0 17 0 0 31 2
1187 188
1158 188
1 4 14 0 0 8320 0 3 22 0 0 5
1132 594
1137 594
1137 500
1074 500
1074 492
4 0 4 0 0 0 0 20 0 0 27 3
1176 91
1176 95
1211 95
0 4 4 0 0 0 0 0 17 26 0 3
1246 220
1211 220
1211 212
0 1 4 0 0 0 0 0 22 26 0 3
1246 296
1074 296
1074 429
0 1 4 0 0 8320 0 0 21 27 0 3
1211 134
1246 134
1246 316
0 1 4 0 0 0 0 0 17 28 0 4
1176 14
1176 24
1211 24
1211 149
1 1 4 0 0 0 0 4 20 0 0 3
1158 14
1176 14
1176 28
6 1 15 0 0 4224 0 17 16 0 0 5
1235 170
1288 170
1288 198
1300 198
1300 190
6 1 16 0 0 4224 0 20 19 0 0 3
1200 49
1297 49
1297 43
0 3 13 0 0 4096 0 0 20 32 0 5
1158 274
1158 149
1141 149
1141 67
1152 67
0 3 13 0 0 4096 0 0 21 34 0 7
1006 465
1006 283
1150 283
1150 274
1158 274
1158 355
1222 355
3 2 17 0 0 8320 0 15 21 0 0 4
1143 260
1166 260
1166 337
1222 337
3 3 13 0 0 20608 0 22 34 0 0 6
1050 468
1006 468
1006 465
979 465
979 530
156 530
6 2 18 0 0 4224 0 24 22 0 0 4
975 458
1021 458
1021 450
1050 450
1 0 8 0 0 0 0 24 0 0 43 3
919 445
894 445
894 253
3 0 19 0 0 8192 0 24 0 0 44 3
919 463
848 463
848 300
9 0 20 0 0 4096 0 36 0 0 52 4
453 286
97 286
97 287
82 287
11 1 7 0 0 0 0 35 25 0 0 5
852 189
954 189
954 103
968 103
968 55
1 2 21 0 0 8320 0 10 36 0 0 4
318 52
440 52
440 223
453 223
3 1 22 0 0 8320 0 36 9 0 0 4
453 232
323 232
323 92
314 92
1 4 23 0 0 4224 0 8 36 0 0 4
316 115
445 115
445 241
453 241
10 1 8 0 0 0 0 35 29 0 0 7
852 198
894 198
894 253
959 253
959 177
971 177
971 169
12 1 19 0 0 12416 0 36 28 0 0 7
517 241
571 241
571 300
965 300
965 236
972 236
972 228
0 2 20 0 0 4224 0 0 30 52 0 4
82 154
567 154
567 224
573 224
1 1 24 0 0 12416 0 1 30 0 0 6
136 129
290 129
290 139
547 139
547 206
573 206
1 4 25 0 0 4224 0 6 35 0 0 4
316 16
679 16
679 180
788 180
5 0 26 0 0 4096 0 36 0 0 49 2
453 250
399 250
1 1 26 0 0 8320 0 7 36 0 0 8
353 370
399 370
399 247
399 247
399 298
399 298
399 214
453 214
2 0 20 0 0 0 0 33 0 0 52 2
210 216
82 216
2 0 20 0 0 0 0 32 0 0 52 2
210 268
82 268
1 2 20 0 0 0 0 11 31 0 0 5
64 122
82 122
82 347
210 347
210 319
3 6 27 0 0 12416 0 33 36 0 0 4
259 207
326 207
326 259
453 259
3 8 28 0 0 12416 0 31 36 0 0 4
259 310
274 310
274 277
453 277
3 7 29 0 0 12416 0 32 36 0 0 4
259 259
326 259
326 268
453 268
1 1 30 0 0 4224 0 12 31 0 0 4
128 321
204 321
204 301
210 301
1 1 31 0 0 4224 0 13 32 0 0 4
130 258
203 258
203 250
210 250
1 1 32 0 0 4224 0 14 33 0 0 4
130 194
192 194
192 198
210 198
25
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
136 167 173 191
146 175 162 191
2 B2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
134 223 171 247
144 231 160 247
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
142 294 179 318
152 302 168 318
2 BO
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
63 95 92 119
73 103 81 119
1 M
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
259 26 296 50
269 34 285 50
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
259 100 296 124
269 108 285 124
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
260 -5 297 19
270 3 286 19
2 A3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
134 100 171 124
144 108 160 124
2 B3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
986 192 1023 216
996 200 1012 216
2 S2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
990 318 1027 342
1000 326 1016 342
2 S0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
972 13 1033 37
982 21 1022 37
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
260 74 297 98
270 82 286 98
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 21
780 3 969 27
790 11 958 27
21 ADDER,SUBTRACT.OUTPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
1312 426 1381 450
1322 434 1370 450
6 Z FLAG
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1317 322 1402 346
1327 330 1391 346
8 OVERFLOW
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 5
1306 36 1367 60
1316 44 1356 60
5 CARRY
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 8
1314 176 1399 200
1324 184 1388 200
8 SIGN BIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
986 246 1023 270
996 254 1012 270
2 S1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
983 121 1020 145
993 129 1009 145
2 S3
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
167 18 276 42
177 26 265 42
11 LOGIC INPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
90 359 199 383
100 367 188 383
11 LOGIC INPUT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
98 563 167 587
108 571 156 587
6 PULSER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
433 298 542 322
443 306 531 322
11 4 BIT ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 11
784 94 893 118
794 102 882 118
11 4 BIT ADDER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 9
34 63 124 86
47 73 110 88
9 CTRL. IP.
0
2048 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
