CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
150 110 30 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 1 0
20 Package,Description,
10 G:\BOM.DAT
0 7
2 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
38
13 Logic Switch~
5 943 158 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V1
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
43332.7 0
0
13 Logic Switch~
5 891 158 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V2
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
43332.7 1
0
13 Logic Switch~
5 831 159 0 1 11
0 12
0
0 0 21360 0
2 0V
-7 -17 7 -9
2 V3
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3124 0 0
2
43332.7 2
0
13 Logic Switch~
5 773 161 0 1 11
0 4
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V4
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
3421 0 0
2
43332.7 3
0
13 Logic Switch~
5 714 162 0 1 11
0 10
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V5
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
8157 0 0
2
43332.7 4
0
13 Logic Switch~
5 652 164 0 1 11
0 9
0
0 0 21360 0
2 0V
-7 -17 7 -9
2 V6
-7 -27 7 -19
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5572 0 0
2
43332.7 5
0
12 Hex Display~
7 1048 508 0 16 19
10 8 7 6 5 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8901 0 0
2
43332.7 6
0
7 Ground~
168 319 202 0 1 3
0 2
0
0 0 53360 0
0
4 GND5
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
7361 0 0
2
43332.7 7
0
12 Hex Display~
7 457 158 0 16 19
10 4 10 9 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-19 -38 16 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
4747 0 0
2
43332.7 8
0
7 Ground~
168 1092 237 0 1 3
0 2
0
0 0 53360 0
0
4 GND4
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
972 0 0
2
43332.7 9
0
12 Hex Display~
7 1040 194 0 16 19
10 3 11 12 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
3472 0 0
2
43332.7 10
0
7 Ground~
168 338 415 0 1 3
0 2
0
0 0 53360 0
0
4 GND3
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
9998 0 0
2
43332.7 11
0
4 4008
219 370 344 0 14 29
0 2 2 2 20 2 2 2 19 16
15 13 30 31 32
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U8
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3536 0 0
2
43332.7 12
0
5 4081~
219 495 487 0 3 22
0 17 18 16
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U7A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 6 0
1 U
4597 0 0
2
43332.7 13
0
5 4030~
219 569 483 0 3 22
0 17 18 5
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2D
26 -6 47 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
3835 0 0
2
43332.7 14
0
14 Logic Display~
6 346 575 0 1 2
10 13
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
43332.7 15
0
14 Logic Display~
6 418 571 0 1 2
10 15
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
43332.7 16
0
5 4081~
219 395 242 0 3 22
0 12 9 19
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U6D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 5 0
1 U
9323 0 0
2
43332.7 17
0
14 Logic Display~
6 598 578 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
317 0 0
2
43332.7 18
0
7 Ground~
168 482 419 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3108 0 0
2
43332.7 19
0
5 4081~
219 473 242 0 3 22
0 10 12 21
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U6B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 5 0
1 U
4299 0 0
2
43332.7 20
0
5 4081~
219 534 243 0 3 22
0 11 9 22
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U6A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 5 0
1 U
9672 0 0
2
43332.7 21
0
4 4008
219 526 344 0 14 29
0 2 2 2 22 2 2 2 21 14
18 20 33 34 35
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U5
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
7876 0 0
2
43332.7 22
0
14 Logic Display~
6 786 579 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
6369 0 0
2
43332.7 23
0
5 4030~
219 762 485 0 3 22
0 24 23 6
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2B
26 -6 47 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
9172 0 0
2
43332.7 24
0
5 4081~
219 687 490 0 3 22
0 23 24 17
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 4 0
1 U
7100 0 0
2
43332.7 25
0
7 Ground~
168 665 422 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 1 0 0 0
3 GND
3820 0 0
2
43332.7 26
0
5 4081~
219 596 243 0 3 22
0 3 9 24
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 4 0
1 U
7678 0 0
2
43332.7 27
0
5 4081~
219 663 244 0 3 22
0 11 10 26
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
961 0 0
2
43332.7 28
0
5 4081~
219 731 244 0 3 22
0 12 4 27
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3178 0 0
2
43332.7 29
0
4 4008
219 707 342 0 14 29
0 2 2 2 27 2 2 2 26 25
23 14 36 37 38
0
0 0 4848 0
4 4008
-14 -60 14 -52
2 U1
-7 -61 7 -53
0
15 DVDD=16;DGND=8;
126 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i %7i %8i %9i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 1 3 5 7 15 2 4 6 9
10 11 12 13 14 1 3 5 7 15
2 4 6 9 10 11 12 13 14 0
65 0 0 512 1 0 0 0
1 U
3409 0 0
2
43332.7 30
0
14 Logic Display~
6 903 576 0 1 2
10 7
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3951 0 0
2
43332.7 31
0
5 4081~
219 818 331 0 3 22
0 28 29 25
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U3D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 3 0
1 U
8885 0 0
2
43332.7 32
0
5 4081~
219 809 243 0 3 22
0 3 10 29
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U3C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 3 0
1 U
3780 0 0
2
43332.7 33
0
5 4081~
219 881 244 0 3 22
0 11 4 28
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U3B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9265 0 0
2
43332.7 34
0
5 4081~
219 951 246 0 3 22
0 3 4 8
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U3A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
9442 0 0
2
43332.7 35
0
5 4030~
219 880 327 0 3 22
0 28 29 7
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U2A
26 -6 47 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
9424 0 0
2
43332.7 36
0
14 Logic Display~
6 968 576 0 1 2
10 8
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9968 0 0
2
43332.7 37
0
75
1 0 3 0 0 8192 0 11 0 0 75 3
1049 218
1049 217
958 217
6 0 2 0 0 4096 0 13 0 0 20 2
338 353
338 356
0 1 4 0 0 8320 0 0 9 62 0 5
722 179
722 173
487 173
487 182
466 182
0 4 5 0 0 4224 0 0 7 23 0 3
572 543
1039 543
1039 532
3 0 6 0 0 8320 0 7 0 0 44 3
1045 532
1045 549
765 549
0 2 7 0 0 4096 0 0 7 64 0 3
883 554
1051 554
1051 532
0 1 8 0 0 8192 0 0 7 73 0 4
967 603
967 604
1057 604
1057 532
4 1 2 0 0 8320 0 9 8 0 0 4
448 182
448 188
319 188
319 196
0 3 9 0 0 4096 0 0 9 31 0 2
454 203
454 182
0 2 10 0 0 8192 0 0 9 41 0 4
507 216
507 190
460 190
460 182
4 1 2 0 0 0 0 11 10 0 0 5
1031 218
1031 253
1072 253
1072 231
1092 231
2 0 11 0 0 8192 0 11 0 0 72 5
1043 218
1043 226
968 226
968 210
908 210
0 3 12 0 0 4096 0 0 11 63 0 5
848 206
1016 206
1016 223
1037 223
1037 218
11 1 13 0 0 8320 0 13 16 0 0 7
402 344
447 344
447 497
325 497
325 600
346 600
346 593
11 9 14 0 0 12416 0 31 23 0 0 6
739 342
743 342
743 400
486 400
486 380
494 380
7 0 2 0 0 0 0 13 0 0 20 4
338 362
338 363
338 363
338 362
5 0 2 0 0 0 0 13 0 0 20 4
338 344
338 345
338 345
338 344
3 0 2 0 0 0 0 13 0 0 20 4
338 326
338 327
338 327
338 326
2 0 2 0 0 0 0 13 0 0 20 4
338 317
338 318
338 318
338 317
1 1 2 0 0 0 0 12 13 0 0 2
338 409
338 308
10 1 15 0 0 8320 0 13 17 0 0 5
402 353
405 353
405 600
418 600
418 589
3 9 16 0 0 12416 0 14 13 0 0 6
493 510
470 510
470 433
330 433
330 380
338 380
3 1 5 0 0 0 0 15 19 0 0 4
572 513
572 604
598 604
598 596
0 1 17 0 0 4224 0 0 14 27 0 3
570 451
502 451
502 465
0 2 18 0 0 4096 0 0 14 26 0 3
563 437
484 437
484 465
10 2 18 0 0 8320 0 23 15 0 0 3
558 353
563 353
563 464
3 1 17 0 0 0 0 26 15 0 0 8
685 513
685 517
618 517
618 451
570 451
570 451
581 451
581 464
3 8 19 0 0 8320 0 18 13 0 0 5
393 265
393 277
289 277
289 371
338 371
11 4 20 0 0 12416 0 23 13 0 0 6
558 344
562 344
562 283
330 283
330 335
338 335
0 1 12 0 0 0 0 0 18 40 0 3
462 208
402 208
402 220
0 2 9 0 0 4224 0 0 18 43 0 3
524 203
384 203
384 220
7 0 2 0 0 0 0 23 0 0 37 2
494 362
482 362
6 0 2 0 0 0 0 23 0 0 37 2
494 353
482 353
5 0 2 0 0 0 0 23 0 0 37 2
494 344
482 344
3 0 2 0 0 0 0 23 0 0 37 4
494 326
477 326
477 327
482 327
2 0 2 0 0 0 0 23 0 0 37 2
494 317
482 317
1 1 2 0 0 0 0 23 20 0 0 3
494 308
482 308
482 413
8 3 21 0 0 8320 0 23 21 0 0 3
494 371
471 371
471 265
3 4 22 0 0 8320 0 22 23 0 0 5
532 266
532 289
486 289
486 335
494 335
0 2 12 0 0 4224 0 0 21 63 0 3
738 208
462 208
462 220
0 1 10 0 0 4224 0 0 21 60 0 3
652 216
480 216
480 220
0 1 11 0 0 8192 0 0 22 61 0 4
671 184
671 187
541 187
541 221
0 2 9 0 0 0 0 0 22 59 0 3
585 203
523 203
523 221
3 1 6 0 0 0 0 25 24 0 0 4
765 515
765 604
786 604
786 597
1 0 23 0 0 8192 0 26 0 0 48 3
694 468
694 454
756 454
2 0 24 0 0 4096 0 26 0 0 47 2
676 468
676 437
3 1 24 0 0 8320 0 28 25 0 0 4
594 266
594 437
774 437
774 466
10 2 23 0 0 8320 0 31 25 0 0 3
739 351
756 351
756 466
3 9 25 0 0 8320 0 33 31 0 0 5
816 354
816 393
668 393
668 378
675 378
7 0 2 0 0 0 0 31 0 0 55 2
675 360
665 360
6 0 2 0 0 0 0 31 0 0 55 4
675 351
677 351
677 351
665 351
5 0 2 0 0 0 0 31 0 0 55 4
675 342
677 342
677 342
665 342
3 0 2 0 0 0 0 31 0 0 55 4
675 324
677 324
677 324
665 324
2 0 2 0 0 0 0 31 0 0 55 4
675 315
677 315
677 315
665 315
1 1 2 0 0 0 0 31 27 0 0 3
675 306
665 306
665 416
3 8 26 0 0 4224 0 29 31 0 0 3
661 267
661 369
675 369
3 4 27 0 0 12416 0 30 31 0 0 5
729 267
729 273
670 273
670 333
675 333
0 1 3 0 0 8320 0 0 28 70 0 4
818 193
818 199
603 199
603 221
1 2 9 0 0 0 0 6 28 0 0 5
664 164
681 164
681 178
585 178
585 221
0 2 10 0 0 0 0 0 29 69 0 4
729 192
729 193
652 193
652 222
0 1 11 0 0 4224 0 0 29 72 0 3
908 184
670 184
670 222
0 2 4 0 0 0 0 0 30 74 0 3
801 179
720 179
720 222
1 1 12 0 0 0 0 3 30 0 0 5
843 159
848 159
848 207
738 207
738 222
3 1 7 0 0 4224 0 37 32 0 0 4
883 357
883 604
903 604
903 594
0 1 28 0 0 4224 0 0 33 68 0 3
879 287
825 287
825 309
0 2 29 0 0 4096 0 0 33 67 0 2
807 274
807 309
2 3 29 0 0 8320 0 37 34 0 0 4
874 308
874 274
807 274
807 266
3 1 28 0 0 0 0 35 37 0 0 4
879 267
879 295
892 295
892 308
1 2 10 0 0 0 0 5 34 0 0 4
726 162
726 192
798 192
798 221
0 1 3 0 0 0 0 0 34 75 0 3
958 193
816 193
816 221
2 0 4 0 0 0 0 35 0 0 74 2
870 222
870 179
1 1 11 0 0 0 0 2 35 0 0 5
903 158
908 158
908 211
888 211
888 222
3 1 8 0 0 4224 0 36 38 0 0 4
949 269
949 603
968 603
968 594
1 2 4 0 0 0 0 4 36 0 0 5
785 161
801 161
801 179
940 179
940 224
1 1 3 0 0 0 0 1 36 0 0 3
955 158
958 158
958 224
21
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
927 104 964 128
937 112 953 128
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
874 102 911 126
884 110 900 126
2 A1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
813 102 850 126
823 110 839 126
2 A2
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
758 102 795 126
768 110 784 126
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
696 105 733 129
706 113 722 129
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
632 106 669 130
642 114 658 130
2 B2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
804 358 895 378
813 365 885 379
12 Half Adder 1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
669 401 758 421
677 408 749 422
12 Full Adder 1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
478 397 567 417
486 405 558 419
12 Full Adder 2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
327 390 418 410
336 397 408 411
12 Full Adder 3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
955 601 984 621
963 609 975 623
2 P0
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
887 604 918 624
896 611 908 625
2 P1
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
774 605 803 625
782 612 794 626
2 P2
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
583 606 614 626
592 614 604 628
2 P3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
331 602 360 622
339 610 351 624
2 P5
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 2
410 604 439 624
418 612 430 626
2 P4
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
458 511 547 531
466 518 538 532
12 Half Adder 3
-11 0 0 0 400 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 12
678 511 767 531
686 518 758 532
12 Half Adder 2
-19 0 0 0 700 0 0 0 0 3 2 1 49
11 Courier New
0 0 0 24
523 626 810 659
534 634 798 655
24 3 BIT MULTIPLIER CIRCUIT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
414 143 437 165
421 150 429 166
1 B
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 1
1027 124 1050 146
1034 131 1042 147
1 A
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
