CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
80 0 3 110 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
0 4 0.500000 0.500000
344 176 457 273
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 805 537 0 1 11
0 3
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V6
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
5130 0 0
2
5.89858e-315 0
0
13 Logic Switch~
5 804 496 0 1 11
0 11
0
0 0 21360 0
2 0V
-6 -16 8 -8
2 V3
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -1 0
1 V
391 0 0
2
5.89858e-315 0
0
13 Logic Switch~
5 800 458 0 10 11
0 12 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V2
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3124 0 0
2
5.89858e-315 0
0
13 Logic Switch~
5 318 159 0 10 11
0 6 0 0 0 0 0 0 0 0
1
0
0 0 21360 0
2 5V
-6 -16 8 -8
2 V4
-6 -26 8 -18
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 1 0 -2 0
1 V
3421 0 0
2
43325.8 0
0
12 Hex Display~
7 325 427 0 18 19
10 4 5 2 3 0 0 0 0 0
0 1 1 0 1 1 0 1 2
0
0 0 53856 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 1 0 0 0
4 DISP
8157 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 749 333 0 1 2
10 18
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L11
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5572 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 748 291 0 1 2
10 10
0
0 0 53856 0
6 100MEG
3 -16 45 -8
3 L10
-10 -21 11 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
8901 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 747 250 0 1 2
10 17
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L9
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
7361 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 746 207 0 1 2
10 16
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L8
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
4747 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 745 165 0 1 2
10 15
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L7
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
972 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 745 124 0 1 2
10 14
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L6
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3472 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 745 79 0 1 2
10 13
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L5
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
9998 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 743 33 0 1 2
10 9
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3536 0 0
2
5.89858e-315 0
0
7 74LS138
19 913 440 0 14 29
0 2 5 4 12 11 3 18 10 17
16 15 14 13 9
0
0 0 5104 0
6 74F138
-21 -61 21 -53
2 U3
-7 -71 7 -63
0
15 DVCC=16;DGND=8;
114 %D [%16bi %8bi %1i %2i %3i %4i %5i %6i]
+ [%16bo %1o %2o %3o %4o %5o %6o %7o %8o %9o %10o %11o %12o %13o %14o] %M
0
12 type:digital
5 DIP16
29

0 3 2 1 6 5 4 7 9 10
11 12 13 14 15 3 2 1 6 5
4 7 9 10 11 12 13 14 15 0
65 0 0 0 1 0 0 0
1 U
4597 0 0
2
5.89858e-315 0
0
14 Logic Display~
6 522 383 0 1 2
10 5
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3835 0 0
2
43325.8 1
0
14 Logic Display~
6 438 380 0 1 2
10 4
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
3670 0 0
2
43325.8 2
0
14 Logic Display~
6 652 376 0 1 2
10 2
0
0 0 53856 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 1 0 0 0
1 L
5616 0 0
2
43325.8 3
0
5 4027~
219 589 251 0 7 32
0 20 6 7 6 21 2 22
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U2A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 2 0
1 U
9323 0 0
2
43325.8 4
0
5 4027~
219 501 252 0 7 32
0 23 6 8 6 24 5 7
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1B
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 7 6 3 5 4 2 1 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 2 1 0
1 U
317 0 0
2
43325.8 5
0
5 4027~
219 422 252 0 7 32
0 25 6 19 6 26 4 8
0
0 0 4720 0
4 4027
7 -60 35 -52
3 U1A
22 -61 43 -53
0
15 DVDD=16;DGND=8;
73 %D [%16bi %8bi %1i %2i %3i %4i %5i][%16bo %1o %2o %3o %4o %5o %6o %7o] %M
0
12 type:digital
5 DIP16
32

0 9 10 13 11 12 14 15 9 10
13 11 12 14 15 7 6 3 5 4
2 1 0 0 0 0 0 0 0 0
0 0 0
65 0 0 512 2 1 1 0
1 U
3108 0 0
2
43325.8 6
0
7 Pulser~
4 317 234 0 10 12
0 27 28 19 29 0 0 5 5 3
8
0
0 0 4656 0
0
2 V1
-7 -28 7 -20
0
0
0
0
0
4 SIP2
9

0 1 2 3 4 1 2 3 4 0
0 0 0 512 1 0 0 0
1 V
4299 0 0
2
43325.8 7
0
30
1 0 2 0 0 8208 0 14 0 0 3 3
881 413
881 400
652 400
0 4 3 0 0 8320 0 0 5 16 0 4
835 537
835 545
316 545
316 451
0 3 2 0 0 8320 0 0 5 7 0 4
652 399
652 474
322 474
322 451
0 1 4 0 0 8192 0 0 5 19 0 4
456 431
456 464
334 464
334 451
0 1 5 0 0 4096 0 0 15 8 0 3
540 410
522 410
522 401
0 1 4 0 0 0 0 0 16 19 0 3
456 406
438 406
438 398
1 6 2 0 0 0 0 17 18 0 0 5
652 394
652 399
627 399
627 233
619 233
0 2 5 0 0 8192 0 0 5 20 0 4
540 409
540 469
328 469
328 451
4 0 6 0 0 8192 0 18 0 0 28 3
565 233
557 233
557 214
4 0 6 0 0 0 0 19 0 0 29 3
477 234
472 234
472 216
0 4 6 0 0 0 0 0 20 27 0 3
390 216
390 234
398 234
7 3 7 0 0 12416 0 19 18 0 0 4
525 216
536 216
536 224
565 224
7 3 8 0 0 12416 0 20 19 0 0 4
446 216
458 216
458 225
477 225
14 1 9 0 0 8320 0 14 13 0 0 5
951 476
1007 476
1007 59
743 59
743 51
1 8 10 0 0 8320 0 7 14 0 0 5
748 309
748 311
969 311
969 422
951 422
1 6 3 0 0 0 0 1 14 0 0 3
817 537
875 537
875 476
1 5 11 0 0 4224 0 2 14 0 0 4
816 496
867 496
867 467
875 467
1 4 12 0 0 4224 0 3 14 0 0 2
812 458
881 458
6 3 4 0 0 12416 0 20 14 0 0 4
452 234
456 234
456 431
881 431
6 2 5 0 0 12416 0 19 14 0 0 6
531 234
541 234
541 409
854 409
854 422
881 422
1 13 13 0 0 12416 0 12 14 0 0 5
745 97
745 109
999 109
999 467
951 467
1 12 14 0 0 12416 0 11 14 0 0 5
745 142
745 149
993 149
993 458
951 458
1 11 15 0 0 12416 0 10 14 0 0 5
745 183
745 191
987 191
987 449
951 449
10 1 16 0 0 12416 0 14 9 0 0 5
951 440
981 440
981 234
746 234
746 225
1 9 17 0 0 8320 0 8 14 0 0 5
747 268
747 274
975 274
975 431
951 431
7 1 18 0 0 12416 0 14 6 0 0 5
951 413
963 413
963 354
749 354
749 351
0 2 6 0 0 4096 0 0 20 29 0 3
390 159
390 216
398 216
0 2 6 0 0 4096 0 0 18 29 0 4
472 159
557 159
557 215
565 215
1 2 6 0 0 4224 0 4 19 0 0 4
330 159
472 159
472 216
477 216
3 3 19 0 0 4224 0 21 20 0 0 2
341 225
398 225
0
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
