CircuitMaker Text
5.6
Probes: 0
41 35 62 4 97 108 86 46 82 16 73 113 113 59 105 107 
0 5 0 1e+09 0.001 2
33
13 10 13 12 18 10 20 20 12 20 
10 13 13 10 20 13 46 20 14 20 
18 17 14 16 20 20 20 20 10 13 
20 18 11 
0 0 30 100 10
176 80 1364 707
7 5.000 V
7 5.000 V
3 GND
0 0
24 100 0 0 0
20 Package,Description,
42 C:\Program Files\CircuitMaker 2000\BOM.DAT
0 7
2 4 0.499203 0.500000
344 176 1532 488
9437202 0
0
6 Title:
5 Name:
0
0
0
21
13 Logic Switch~
5 543 168 0 1 11
0 7
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V4
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
9840 0 0
2
43340.7 0
0
13 Logic Switch~
5 597 165 0 1 11
0 8
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V3
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
6910 0 0
2
43340.7 0
0
13 Logic Switch~
5 661 164 0 1 11
0 9
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V2
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
449 0 0
2
43340.7 0
0
13 Logic Switch~
5 725 165 0 1 11
0 10
0
0 0 21360 270
2 0V
-6 -21 8 -13
2 V1
-6 -31 8 -23
0
0
25 *0=0V 1=5V
%D %1 0 DC %V
0
0
0
3

0 1 1 0
86 0 0 0 0 0 -1 0
1 V
8761 0 0
2
43340.7 0
0
7 Ground~
168 686 108 0 1 3
0 2
0
0 0 53360 0
0
4 GND2
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
6748 0 0
2
43340.7 0
0
7 Ground~
168 561 112 0 1 3
0 2
0
0 0 53360 0
0
4 GND1
-14 -26 14 -18
0
4 GND;
0
0
0
0
3

0 1 1 0
0 0 0 0 0 0 0 0
3 GND
7393 0 0
2
43340.7 0
0
12 Hex Display~
7 569 74 0 16 19
10 8 7 2 15 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP3
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 512 0 0 0 0
4 DISP
7699 0 0
2
43340.7 0
0
12 Hex Display~
7 691 72 0 16 19
10 10 9 2 2 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP2
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
6638 0 0
2
43340.7 0
0
12 Hex Display~
7 820 316 0 16 19
10 6 5 4 3 0 0 0 0 0
0 1 1 1 1 1 1
0
0 0 53872 0
4 1MEG
-15 -42 13 -34
5 DISP1
-18 -38 17 -30
0
0
50 %DA %1 0 %V
%DB %2 0 %V
%DC %3 0 %V
%DD %4 0 %V
0
0
0
9

0 1 2 3 4 1 2 3 4 0
82 0 0 0 0 0 0 0
4 DISP
4595 0 0
2
43340.7 0
0
5 4030~
219 507 309 0 3 22
0 12 11 4
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U3B
26 -6 47 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 3 0
1 U
9395 0 0
2
43340.7 0
0
5 4081~
219 441 314 0 3 22
0 12 11 3
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 4 0
1 U
3303 0 0
2
43340.7 0
0
14 Logic Display~
6 459 401 0 1 2
10 3
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L4
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
4498 0 0
2
43340.7 0
0
14 Logic Display~
6 531 399 0 1 2
10 4
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L3
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
9728 0 0
2
43340.7 0
0
14 Logic Display~
6 666 396 0 1 2
10 5
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L2
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3789 0 0
2
43340.7 0
0
5 4081~
219 580 308 0 3 22
0 14 13 12
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U4A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 4 0
1 U
3978 0 0
2
43340.7 0
0
5 4030~
219 646 302 0 3 22
0 14 13 5
0
0 0 624 270
4 4030
-7 -24 21 -16
3 U3A
26 -6 47 2
0
15 DVDD=14;DGND=7;
49 %D [%14bi %7bi %1i %2i]
+ [%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 3 0
1 U
3494 0 0
2
43340.7 0
0
14 Logic Display~
6 758 395 0 1 2
10 6
0
0 0 53872 0
6 100MEG
3 -16 45 -8
2 L1
-7 -21 7 -13
0
0
10 %D %1 0 %V
0
0
0
3

0 1 1 0
82 0 0 0 0 0 0 0
1 L
3507 0 0
2
43340.7 0
0
5 4081~
219 482 236 0 3 22
0 9 7 11
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U2D
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 12 13 11 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 4 2 0
1 U
5151 0 0
2
43340.7 0
0
5 4081~
219 579 234 0 3 22
0 10 7 13
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U2C
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 8 9 10 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 3 2 0
1 U
3701 0 0
2
43340.7 0
0
5 4081~
219 664 233 0 3 22
0 9 8 14
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U2B
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 5 6 4 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 2 2 0
1 U
8585 0 0
2
43340.7 0
0
5 4081~
219 742 228 0 3 22
0 10 8 6
0
0 0 624 270
4 4081
-7 -24 21 -16
3 U2A
16 -4 37 4
0
15 DVDD=14;DGND=7;
45 %D [%14bi %7bi %1i %2i][%14bo %1o %2o %3o] %M
0
12 type:digital
5 DIP14
22

0 1 2 3 1 2 3 5 6 4
8 9 10 12 13 11 0 0 0 0
0 1 0
65 0 0 0 4 1 2 0
1 U
8809 0 0
2
43340.7 0
0
31
4 1 3 0 0 8320 0 9 12 0 0 4
811 340
811 437
459 437
459 419
3 0 4 0 0 8320 0 9 0 0 13 4
817 340
817 432
531 432
531 425
2 0 5 0 0 8320 0 9 0 0 14 4
823 340
823 428
664 428
664 423
1 0 6 0 0 4096 0 9 0 0 15 4
829 340
829 418
757 418
757 421
1 4 2 0 0 4096 0 5 8 0 0 3
686 102
686 96
682 96
1 3 2 0 0 0 0 5 8 0 0 3
686 102
686 96
688 96
1 3 2 0 0 4224 0 6 7 0 0 3
561 106
561 98
566 98
1 2 7 0 0 12416 0 1 7 0 0 4
543 180
543 189
572 189
572 98
1 1 8 0 0 4096 0 7 2 0 0 4
578 98
578 190
597 190
597 177
0 2 9 0 0 12288 0 0 8 24 0 4
661 185
661 180
694 180
694 96
1 1 10 0 0 12288 0 4 8 0 0 4
725 177
725 181
700 181
700 96
1 3 3 0 0 0 0 12 11 0 0 4
459 419
459 421
439 421
439 337
3 1 4 0 0 0 0 10 13 0 0 4
510 339
510 425
531 425
531 417
3 1 5 0 0 0 0 16 14 0 0 4
649 332
649 423
666 423
666 414
3 1 6 0 0 4224 0 21 17 0 0 4
740 251
740 421
758 421
758 413
0 2 11 0 0 4224 0 0 11 18 0 3
480 269
430 269
430 292
0 1 12 0 0 8320 0 0 11 19 0 4
521 277
521 281
448 281
448 292
3 2 11 0 0 0 0 18 10 0 0 4
480 259
480 277
501 277
501 290
3 1 12 0 0 0 0 15 10 0 0 6
578 331
578 338
535 338
535 277
519 277
519 290
0 2 13 0 0 8192 0 0 15 21 0 3
577 265
569 265
569 286
3 2 13 0 0 8320 0 19 16 0 0 4
577 257
577 265
640 265
640 283
0 1 14 0 0 4224 0 0 15 23 0 3
662 270
587 270
587 286
3 1 14 0 0 0 0 20 16 0 0 4
662 256
662 270
658 270
658 283
0 1 9 0 0 4224 0 0 18 29 0 3
661 185
489 185
489 214
0 2 7 0 0 0 0 0 18 26 0 3
543 204
471 204
471 214
1 2 7 0 0 0 0 1 19 0 0 4
543 180
543 204
568 204
568 212
0 1 10 0 0 4224 0 0 19 31 0 3
725 197
586 197
586 212
0 2 8 0 0 0 0 0 20 30 0 2
653 193
653 211
1 1 9 0 0 0 0 3 20 0 0 4
661 176
661 203
671 203
671 211
1 2 8 0 0 8320 0 2 21 0 0 4
597 177
597 193
731 193
731 206
1 1 10 0 0 0 0 4 21 0 0 4
725 177
725 198
749 198
749 206
6
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 6
784 249 853 273
794 257 842 273
6 RESULT
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 16
562 455 711 479
572 463 700 479
16 2 BIT MULTIPLIER
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
577 96 614 120
587 104 603 120
2 B0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
525 96 562 120
535 104 551 120
2 B1
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
706 97 743 121
716 105 732 121
2 A0
16 8 0 0 0 0 0 0 0 0 0 0 54
11 Courier New
0 0 0 2
644 94 681 118
654 102 670 118
2 A1
0
2049 0 0
0
0
0
0 0 0
0
0 0 0
0 0 0 0
0 0 0 0
0
0
0 0 0
0 0 0
0
0
0 0 0 0
0
0 0 0 0 0
0 0 0 0
0
0 0 0
0
0 0 0
0 0 0 0 0 0 0 0 0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
0 0 0 0 0 0
0 0 0 0
0 0 0 0
0 0
0 0
0 0
0 0
0 0
0 0 0 0 0 0
0 0
0 0 0
0
